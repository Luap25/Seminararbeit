PK   �-Z����  R�     cirkitFile.jsonŝm��6���B�rX��&����p�]�E�v��,Q]]��+�yi������.ۼ�5�tW�R�Ù�HV>GM��-�q��]���Et��$zʚ�C�4�D�j��֏�5��)�����OK���^�E�h$��Y��NcY�:�ti�(�Js���It{�n�����q��.q�
����5N���-,vH�<�$�!�cH�>���!�cH�8�?��{H�8�?��#��H���oT�P�扈�ճX3�<���0\����ӏ��`�֨�-�k��Z$�Gu�0]KT��u����r���%.�!F C�@��1b$2�Hlr��O"��H�$�?��O"�S�s^g<_��Dt}��*D�g�}`xFt}a���9̤��!]_X�!�jXF��ds��x����L�+��&:H�B�	�Gi����Dc�0��/D� }$���e[���y� ��7I��P�H+�Ċ �"I�(+)�MbŐX�4��KC/������h f43�ÌbFC1����`�9Ŝ�bNC1���w[�$"Ø�(.K+�Ø�(��H�&��RX���b��Ę���8�p��ł�bAC���ł�_,i|���Œ�K����bIC���X�P,i(�4��V"�����╸X��K}�"������X����RޕL"�*G0��K �FGa�#��Q���7`kZƣ0�^͆Cs����`k��֭ڬu�j�­�&�#�ux+�Ċ �"I�(+)�MbŐX�4��KC/������h f43�ÌbFC1����`�9Ŝ�bNC1����P�i(�4�ł(���X�P,h(4�ł�bIC���X�P,�2b�%Œ�bIC���X�P��SZ��[��B�ux+�Bh�o��2���\_��:���K �ZG`��ހ�ap����[��j�����պ���	���ퟬ{���ѭ�D�ƭ��,w�c�x���5��=�y��3��$�.�Bg��E[�]�f��l��<��7\PO�y�
�5��k��}y���Lx��'<��c��]A��� ��q��VPg��������5�~�.[cN���y�w�w���`H?��v#�>�:��W�w�0��/�G ��9P���v_e5�Fǯ�C���[����`ȐIp���`�ԇЬ)��b{��{]���Q�uU`xD>���H}�ԗH}��O���o���@,�� �2Ȱ2,��!�rȰ 2,�K"G�B,�K"ǒȱ$r,��m������ͩ=L���x?��ʞ�S{�ҟ�[�G��ߠ9��ڳaX��q�e\`���z[����m%��J�����K�Ē(�$J,�K�Ē�.�z�<����9�硷��M�t�d���z;3�K���BLB�c�si-�?G�䕃`	���C�2�����7�Q�r9l�^&�N�*|�
,�|�*�U���x��ݡ��Ҽ���,�?���k����:A/ɼ(��3/ͼ8���+0����l{�5���^�{���ڕ7��^W��j�]�Yx�5��^Cx�5�o-J�!����;�!����kH�!���ކVd��K]�*�E,���MZ�8MJfE2���
�_s�+����]��_��~`'�v:�m�� �{a����Zǽ�
y��4���φ�~�-�^����~�J�^7��I�[j��h���ܯ�ӥ�����)�];m�C?mC�8m�C�<mRC��a ��g�ˊY�5����~�W����[����>k38��;t��K״���M�^Um�/-�K��¤:M��=I%�J�L�X�s����ɢ��б��ؼ��LsJ��3g���/��AM"bm��{CA�l�MV�~��z�mWM>wÙ�˧j���^&z��/�����NᤸT�yʉ�r�SJ�733~Z���)�G'��RI:U�J�����TH?�ͥ�(*�1څ5]�:>nz=k��JٷC��q��k�7?�.��a�ǒnj�]�ڝ�Lu/fƛ��"L­���(6���Slǥxo$�������Rr\Jy[BۤK���t#5n+Mx/�/��2"%�����=�q)9��R$%�\��@�R�o��δ�^_߬4� ��sb�����i����s�S뚥�p=:a�b'�?.vr)��N�;�l\L�\����N��M7+.=#^sa�3b��,��vi��v}E_�c_5.'E���bgXoH��e�{���Q�.r��������|~�ٳ{�n���͟��CT�f��p������il�� +kt�! �N�}\���5�j��{]c�<e�D�vI1��<��p���������W��gE�����VI���d�v��z�\�{ʖτ+�$�Y��R�<6F�q�\V�4�D&�\�^�켉aN@���+�w&���y�g��x�*��\YH(��L6V2e��3:=��WY��훥[�[Im� ��U�!U!�Y.�ب\����l8�C+�����fV
��E�3���E;��8Msn�,3g�p�?|\f��y��Y�Sa���v��c��,o�p�l�����O#?Teՙ�W�i��~�]ݴ�(�ƭVC�˄M$W����Ԧ�t�[�%��.f���2��/ә�EQ*��nv7���O�"�af UW��Yf]��,S7�c�r�� '`jgel���JI�Y)�⦄M��$yʡS�x3..u�$yɎ�/���>D�몸Y�v����o>?<,nn������T�����K�<��Mn���Y/njHxoA�{���������Z��i��e�+����#��.o;��Q�L�I��������X�?x9�Cp�}H��ڷ��m��)$� ��>"zU??C�����^�M��F�~�HL���|��� �&� ������'�T�f�����Ը?�U�~yt��y�T�.�����z�;����S������\룎&Q9���6��*��j��}SͲ��ߚz�(^m�=j7�c��L|Sv��'�S����3�d#��]4����Ǿk�u��Q���}[��F�n�F�]�v����^�"� ��܇K�;��2��Nuj�EN��	d�S��`g��D�a_���3H!v�d�E�)+�L�~�'��.�킃J��w�_�p�g@�ib� �m.Ej���,�)��m�Uy�)�b�X�t��,:�
l���j=�%SۏO����D�l�;�-@��h�Ʀ<��P_�d`7������H5��&��T�rv�(�v%�&܌ڔԃՄ�x7���ʏBqmr
I�:h�����R�H�O�]G�I%B&�`sc7�T+}dBL�2p��C��l+�q!�~�cRù�	̤2�m����j��v����۸�tc�7��֚=�k��R���]�j�e�~{����һ�~YG�[9E��,�K�8��ߞ� ����o-���#�O����,r�w�J�]����/����揯�~�9��.�^ �vX-��Ő�|�m�>#[�m��L5ه��c�?�oYW������C�K�o�;��KNV����{W)�?���o/0�@a�D���V��8��޽@f8�ѿՓ��F�FB��@cW�ڿ���C6���A�����I�"Կ��!�	J�G�P�Em
����%L������������HK
���CS�aH��h�*����HJi5��CO�T��^�.'R��I3i�bt I� �H�j�c�$�����:+u&�t�'�-�N�[,)�·P���^�4���R=~;V��o���5U6�]��e��R����:�W?�nݳ�T߿�D-���.o�w����CI z�PK   �-Z����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   ��-Zl��B�  +   images/60459fb9-c9d0-40e2-ae43-752ef2ed40d9��gTSm.��H����ޤDE��;Q��C�  �	(-*M�Dz'ҥK�^B�	5@��;�?�ǽw��V�z���g��3ϓ�?�ඎ�������� ����������_'��nPP�_��AI�ߛ����������������QRߢ��y���m��^W�M*J�������@EVJ�DN���@F�@F�  ��d�� ��Ȯ�S\�q��5���''�v�u
���Ыu �u�{R�o0����f�~�����IE���_��'�����;��}�B²r�
�J՟>�����16153���rptrvy������!"2�ctLJ꧴��_2����(�YYU]S[W���������otl|br�����
zum}csk{xt|rz�;�������#.�+\׮΀��?\d�������=���)_y3�J��b~������O��b�3B��/�,����D��X��/d����5�INvux� �B��u�/�!��J���0��<��p��I(�Vu%����ɉ�ec0a��l��h	 �I;��t���e�\Aq߂+b&?�[��F�վr`��7O&�T������1�,��X�!n7?�j���[8���<�����^W�3�a�P�98۠�_5Z7�j��2�L.�^�yo�`JO�?']+<=���{,o'�!�e�m�ɵФ%�y��]L���h�'���]��m��h9���Mq�5ٛ����m3I 6Cx��d�y���C����th`��'BNVx�vK�^�Hv.�c��<$>� U��K��M���'�q��Pw �#��\|���	a�t��繹�KV'[�#}�@v���9���k>�����Gp���M�	z��� ������ʤ��ܻ��#.�U_Ӹ�������(�m!|����&v���]�8!�gB9-��q���e.:��,H�Ƴ��Y�{��

)���dܝ.��`�U8x�b�[Hj�9_����<<�N�*�f�%�5>\��(���$���-��{�*�����T��[��
�)���4e0mⲑ)�T��VX�G� 3�����筜M�{A�#v{¿#jߎ����"�)�����7�#P�tk��h�����#�O҂��W���C��svG<�?��طD�0��OW�o�j��������{�fr�~f1�>ܿӓSl+��� н{Ʈsi~ZH(A�� 3�e�����r��6���vI������{����Ͻ�f��Wb@�Z����w�ƒo�o,�`���y�UZD����5��.�n)a�RÒw���裪�x�`NMB2_I�����a���˅N���3Uǲ1��{�� ��@Bf�~?x�c���A������� ���F)T����WV�wc�s���#]�px�z�-���lJ�Ah�DK�pX?��\��q�{��d�tQ<��٩}߷R��E�����r�ij�z�E)���8>n`�F�ϭ����bx�e����إ素H�W2oh��ٿ9 �r��uGH�_e���R���5��M�@�9�T��U���<vQŤ���!:s��4�V�2/ 5`����Q����Q�66���F\71 �,_>���!&�xӼ����jR|gU�Bsƫ��l��3���Y�:��_��E.���{>,�~)��A��oi�^mɀ���U��Xks��JӇ�j*�3����K>/��h������>������
���,��Z�WaQ�����	���Ƒ��4����bPq�r�_�%�Z�ϸ����r�x�0��Fυ�	1�S��Q�b��E���8�{u�E5L�����C���ŵm�Pjd>��hSW�rY�BE�Ć5�$��y۸5:��7�lY��?8���e~&��D0����mpiX��'ѹ��5uI �Cw�ݣw���Qw_���D���Z�h�h?�T��-y}���� �H@��m`l��n/�v����ك"H%��{�_�;����b� AȬ0�&Y~������oP��Eߑ����ldtd�ԭ�����`�o���qϢ00��7���d����+�H��֘f*���d�$�\DP����I�E�k�~��G����N�j�����K�:��!�)D�=�)\o匪d�_��1#�����e.�Dah0�Ŷ��a�� ��'���� �s�4���@߹�(ǀ��χ"������[_�A���4�#��Y�?�L�"p�U����{���@�A�����G׏H_O� �����^��^�iR.�To�����v0-(/=�V�S��?��u��As��Ĝ��nO�2OT#@�*uԜ^����5_���o�]�e������W�E�mJM%آóiF^|k���j�j�R�N?��aC� ¯PI���$�ʄi jU�߷��*O{7�vPO٢yl=!H|�.�h�瀥�~[b�]��:?������utP�1[�B���I��
l^ T�[TtN��m����>�S*��ַ>��<��h��p!o���U�T��)CmB(�ޡ��
=^�v+��� ��#L��e�e�]!��F�����É��o{�H���3s!����o�k��6o9vަ�#����Ԋ�\'����^�m���2&�s�X�Sihܮ�7�;ĩ�w0x̍�n\�:�E��HNA���u�qazu���O=�M����ϓ b�x�_2�\Gt�G��K�v��p���d;c�u�+%�:V�^�Q������
�
���[��ssG�
�<s�e[�M�7Y���D�N�u;��BT��,C��I���>�2��{U�*���\x���xo� �EL� ���u*��9:�����*U{鿇���g�����+��I���I��:��m�|=xO�l��4(�[|H�yʓje�sg�6�6,ۯ�mEy^�`��>)3s�����S[rQ���X�E��=-.E�B�r��r	4p�^�G1�4߈\V�tsHR�����3�7��(Rkpۑ ���j��rD��G>5)N�n?��`�>�#r��ړt���pM�<zy3�eA��j�����L�o��ŭ7#�x��s����~axD��_�ۘ��ړ���%?O4�؀A�_�N�%ųU� �P�K��g�j8SЌw�z�ҭ����ӽ��'�`���w�<�mu��2��!���D���R�<*���($a����1�$ "���kI�+v���ky�kk��뚴��B��i��Ns^��/t��Q����+�=�[|N�B��M�WA)S�
��R�/V�K�A�'�7���2[��|rܡ"-	j�Ս�Zp� Eڔ��!�!����`�u���������|��>"R�{�O��KB��	iY�6G�|9=�\�#�8�e�r�4�9�Ȋ���0UO+������Px���aڶg�J��H`�uB`'�����0��D��4����₱��4���j��~�� c�.�s����4H���'���6�O�Ns��ݛۃ�r��%�tx,{6��x�
�lm�杀���%i����ita3G|VpH��n���.��o�bt�p����/?e]w��/n���-b%�kg�cU`�����SX�5y��'Zo�Xxuz��}\cY�2�K%Y��W�����$m
���$Fd��X�[�ըNd{e�8L�
���r����]��ާ��y�i�"@Nw25���C�D��ҥN%�c�V�3ti��V`Q�%��f���G�=�oō�8=��OW��f]���]I 
��"��$�i�4	9d����=Af��^�U[��Э���$���>.���n������<���p��';�a7-�p�D��	�U�?O�s��8<�Z��g�H�؋��g�;�,EE�ʉ�@T�׵�c�~x�S�� '���� r�:�<0Q��W�J��z7a�{����z�	��XOw����e��|��+�
1yj��M��x�r�gN��tTlyӓ9�KoMPd@!�
�^��D�O0�Yյr}�O!��A�|��ސ�ګ?���w( �^�o\ҢX�M����L�N���	���N���Pw<�P��CI��Wl܇�R�3���p\T�q��<b	�f՚Wb���ݜ����J~�U�x�Ԍ�˴;3�=13��X]֧��ZPM"YWg�/��u`�6�c+����P�d̯ r�;�u��۶\�{|E�Xq���̤:l:�y������3��]z�����ry�
m�ȏ�<21�ʋJ
�,�e�۫QS�ѷ��r�����\��[���u�Ggq*�y����)m{�<������"�9����")ѩe�����O�z׍�*�a��i2Gc=�y�N!���%��Fq]ZSBj� �V����{��:�P�Y�I��H6�gx�Du~)�/�]D�����Lk�E4�e�o8��{�����g�UW����J #�0�_�������켡����ߤ�+�y&#jks��A�:�Gކ�����v���i�0
����	ѵ�w6n���[*�ӵb��+��~�J����Zmw��W���2��?��|�����~��W Kض����})5z�N�I��-��0O��#,+!_c�"D�w�1�tu
ߩl̎h�䶮��HF�Y�0ų��Ǘn��5��WE����Bp#�A��|����R������,�07�������mT��I�T��P#qەcQ`a9��?̣�R�����x���)T�Io�1��Ѯʪ��(]>TZ�i��=ފ�,"R�,7Y����E��ˀ*}��Y��_<D��m�-v��6���yI��&.��������f�6�� �e��Z�Hu�ĩw���u�m���d����=n���zW��C`t�lA|�M+����]�42��o׾L��c�m�0ʀˈ£�X�:�ٻ��|�&�M��\Aj�X��@t��y�����S}K���;�2/}=��q96nUs�4ن�l}.'�C����>�'�_�Pv����!����*��3��vR�G�hο ��Њ;��� O�]�壽0�����{QsT.�kȬU{~O{�Yv��h��#����6k��s��v�;����v,+�+�q����Vi�����u�x����f }a�����#M�\�&�d�wB�uL&e�b
������Je��>}�\�����)�/���_"�U����9�B��87y�Ǘƶ%gw�$�K��m�z�9���d=�?y� |]������wal�W����@�"���u���_$@����>B.J+?����	$��'��i�\��mq�g<x��t���&�A���ˊ����c�p��`��RW��d��[`�aף�^�)�����S`�[+BWKz�ܒ����ˏgs����
��_����V�i�Xs���,#:/�H_�B����MV�ۙ���ޝVݳ�����h;�"h�K�{��1޺�;�,�����;?[YFƴ�v�5׬�ړ���V ��9%_��NV7����f�)����fE���[ǋE��p|�;Cٟ+5�bm�W��_Hy/a����i$L�����h�w�{�����1�����a3��%��z.�{�XQ�L�Y�xC��.����v�?gؖL�PR��}��ˀ2�r��3s�K��2i,�^�M]i�W�mv�����N}���F��mu[#�{[a
]Dc?��/&hJV3�B�C�>�(h~��dxҸ^�#�"Դ�n���H��������C�L�����z`�ܨ��?#D��F��`�6W�7�E��7�kO=�~���3�t��	�j���tp\A�|n���G\@9g�l{���g�'Cw�7��&�m���m+h���Nc�D^����Y6������se����쨃(���жKZ�ޕ��c��2ݏ�&?ϓw��t�qS]AH�|�B(��E�b�Q��v�C3�9�����2��ĕh�]`��_z�^_=��ݎX3��W"@/d�@����$�3=�>��l1�$��C�}7���3�C�Pq���Z�;]�ϯKߪ��6�ϔɏ��p6����7:�T��f��5��%�j�_�c�6���¨�)�Un,��c���Fs�&�����rO�����* �P�\i7��Jaw����ðer)#ybk�S��ܗ:ux��ƨs0���cw���F��'�ݔVM�NxZ��
=N��#1��a��=��Ɩ�}}���7��ˁJ\��wW����c�T��ߛl�\=���k�N��cv��GO�?������׹�G;�y�ņ�XE���
sP,]��M�|@N����Wdy'���*�F�M�kAS��8.��͸�5�>;u���u�Z�ӜP�G?��%h�9�������e�)y����[M5^`̋E��/��xLY�w	q���D���G�z?�0/z���)>�N8`OÚGw�lC��Ls�s�m��R��4�f/���&lė8�#_3���x�(ϭ��o�u�]��kBHsw:"���&ܾ�g�䔷�R�7�Xk���=�,Å���y��� _ɦ=���~pMcse�gZ��_(*~��a��R��&�5p<���Ԟ�
g�gl9�ׯm�@trm��E�%���Lb~`�&�:�Bū�����j���B���T��ѡW4��:�wH�z�����<����Y���M�w�L�(	)�+���ՠ�j�����x�AﳿB07#QG��3�tj�+c͏�p�`��1މ�����*�b�3��\c(��WrH܃��ASq	�\8�+�J��u#7U��g���� ��3�t�99L��ӣ���n��t��
ň|��Y�{`��Т��ț8z���-V-�Pi�<k7���Ɠ�z-�{�{mF핿1����gN����T������H�,�W�z˨��_�V�u�ܰ���O����!�Z5ڢ��)��e�ʑV0�?�c}s���1��\�O���Ș�v�0���
Y4G}<Aƌ�lX6!��ᄟrz�G�?�J(�$���Oϐ_U�t��T\/:�ɳ�-�y4c��[!^E�j��s����C��.�����M�z�N^�j���u�::e �����Akx]�e�ƑQ]0����]Ӥg:���Y�ND6!�0�+��9ie�<\du�d�ѯY��!���Hd�&�d�(Fϲ���y����6��d��[@_h��`|���*�p\D~_ϥoG]̟�逨�R���&�t~�?H6�߲��B %��0v>D.�i�v��4�P�PwEr�Dg��������Ps�^c�+��f 6��n��f+��'>��b��O�Ԉ��%,��P1��>Ԣ��2���e�����zDl���7�YU1�2�����`�N{'A.$ �`Y���%�Yʨ5Xm�O�+��r������*J�e���,���t������ʪ�{"Va�(O���
��)���n���Q����5i�,��k���
�<��y�)�OOu�Q5���9ur@ko�l�>^/Y�\WmxC����D佪�_x�|�Aϻ�s���'?�n����/��A��=�TV��-c�/�%}���%�ԅ�6�����#�
$�ĕf�ezP=^Jl͐ ��v�xtc!�pӿ�>)����H�论� �p�@/��qKXF$u�:zP$,����vW1!�OpK�Hڠ��������r�9���nݕ
��Bf�����Zs��ʍ4�����^�$ɷ�����y�����Eǌ�#�SĤ���n�g�u�e3|3ý��[��VD7F#n��TNѪ�\��=\l���9_B��12���DH���L�e��-��[%NJb��VzM��/C�Q��j®d������z���+���r������Uj���2�=���3$�WW@B�A�x�ŕ�$�nK��Sв�:��yƂ��`'�<��n���@z��6��"��!���Gw���\�MNQ~����n��s�3�����^��~�Dt�3��3�(���D~�5§
��]Φǿë���9�gW�+%��=�|���uWΥ�����/�e���4�⦿���	�$ �T/nK��ݠ�AT�&��>g��F8�/�2��i(�������l�qk_��^q�
���CՂ�]I�Z]��.�ĵ^�Z"����|�w��{	iQ�$ ϖ� ©z�M�y��݆�.S��wt�Pc� �m�5!���o�X"?G*�~i�Sݾ��{�k�X��U���F�)�Ŭ������J	����]Y���*&@�H }gI(S��~:�P��k䪳=c��j��R���9����fm��������/�Mni��ϡ_m������]"��g�.f9W�Uzf�q�$}{�����*�E��+���Oό/p�
썄1�`-�8�9X�ߧ���N���t��?��>_	[[�Ye���)B��u®J�,��fr�΂�N[yeM�����m����X�����;<�m�KG-��h�4C ?���}XP��U�X��+VS�6V������qD~��l_��7X���Dt��~���g~t���ϥT+Dɣ<��$��r)��a�H����:Q��C.�kJs���ME��^����)�K6�`�Ʊ��2�J��Q)����ЭK`??���[7H�s�����
0ߗ�ծS��V���O��qk�Tk�'Y������"g�!	e�0�SO&���?���2q����¤����X��f��o�<�5���N=��-t	Y޾����]�����,���.�AǷՍw�w�o�0ޝ�iD?�7q���7�p�M��7����A�dO����r��V��פ,����IvcN���Q��|֭��]�Z�.B*�3����.*���8ރi5U�j�S�]�AY�P��7�Y������_w���O���+�[��wsZ�7��K�۴���ּ߂h_�n�V�ԍ��]8Pr���g��-200~&�W��J�r��N�v�z��ͻ�ox�wL�˟�U���E/�XGd���q�e��<��Y�AiؖQ������V�\����ؽ1�D���/ĕ\��	9=��r1V�.�Ne�y�qKq2
GJ��nP��N�U���	�[����5z�W;���.����uu��2�NCUˬ�=�'ԩ�n�"n��ɝ�B�����ū�<�#D�E�i����K �WD@B-K��t��rŲZO��N?�����8������6	R��ہ�&~��^Kj��^%[y75]��晊�w�3�t��h� �_���x��͇r-'m�|m�5(�s��k�|�FR5ݏUb}�����:���C��S��.�m�lxM���.���(<C�iԔ�[�jy,{��"��� m��I��,�KW��?j�����E�YG�xiQ=���������*�*�oxӟr�u]�l���>D.�N6U�I�v������E��� �3��c��;�;P�˗���4*�B�(U�N�:�"2Fg� e�ˆ�$�nǋ"����+*!oc���X��p���nA���V�S�6T2��rH�ب��*�]��UL9�%'%q�a����<�
��i�)���/!Ԭ�x�谦�$7�g&���{L�� �ǅ�F����&/�5$��˧GX{�<ܙ�+n36q�Ɇҳ�oS�]_�0Ѯ�k+�6�(fxGL����=�����{K����:�l�Y�1p�{4J���!�1(ʽ�����wbH ��Zזp?w���Ü~��g[ �Y��$�;ԑt�������g���74�i��L�� ����D<C�
��0����VL ��&�\CCK�Dk�cݑn�U���7#��m%��E٬�Hx����G���!�8��=K�A<���w��&����{Gzo.Zf��S��>��(���z_Q�a��\�!��CTm�����'NЎ��_Jl4��r�xCG�A�/�%-�����a�����Ր�Ƌ�K<�,9�u�^����r�4\OqL1���"�"5��2�F�ɝ������c1B�3zVj>����@M����F��Z��+�����#����R��.?$WR�:���w�$�y���}=?���a\��({�=��HC�	\��[U�$����eM�`r���3��mr��Rcɷ��+���|Vu�}Z�6TZ8H��8ܾ���EÖ-(��T���~Q�\����ǘD�{�˓ 4Hj�"Qj�ntJ��jmm�LQ4�vΝs�䁖3���{0`.X8"Q?��Wt���C���:A{	��&Ҹ��W��k G�7F��Ԧ/L��GH �-cQGh+���d�	�XT�Q)�c#����䫁0��&�D;��d0<��y|��{�9��X��nj�[|̴D���3NϫG7/o�5����I�a
�TdFY�p&�6o��r#6Y�����p���/���rXȠ"]
q j]i��%�p�s��:����{v��{*�&���w��|��2Y"�=!E���rvo=�_�'��
<��ˡ��P�B2$m݄C��@��*]  � E�w������(˒c�_�n�kN�Ѵ�c�b���5О�Z��w{b;ܞ^Iw����
X���`0�s��M���w�/{
��P�Ɇ-5QKˆK�p�{�)Jo`�;�V�9bWcP�2cy��%es�=�<	��s�Z����>-	�	�.v��ѽ��ti��T���8�1���59��ۇ��&I�LGY`��4��o�����]"��O9Svޔ���ի}����Lmg��{~"��x$�U�������]�X@������f#b�����֎3~aR�l�@C�w���G�������Y�����2U@'.��>��j��=/*~���5����D�'��(�*V�E7H�T�P!�_��$��*���}�і�:p���H7>�}'$=k%KD�����җ0hn8y�	R�>~�<�J��C�(�R�d��Z�O$��(,���7�0�jCY�+fi���|`��>Ba�+��V�^�6�"fie��V.������>�FЧʄ�wz���?���2*�/��|\������=�2��^�,|J!�b�������TE(d�����ޒM��̿�l��<՟U�dIP�flW�[ٱ�a^q��j2;خ(/�A��V�4��s5$T@������W����4��2�K	ؔ���$�p� lZ��������z����S����Bl�����z�%����b�1=�4pɟ.�)E1<5��ۄ�[�d/k|�K�}��U�*�y��$
��k�I�l��4����c�m�����_���!����-������Hq/@�� L��p����fC��������t�W�e��oЅ��'�����'UAwMS�1�=
�*�;���םpGD�D�)ӌ�|m�+a~WO{��̺�%֏�U?1
j�1���8����H>ơ���A�z}�+.����ֱV.���]�V>@o>�M�����YZ?U�m��9��<�L�3ɁX g�/������]�?�ݥ��(�Ay$�U,C�����[X���=�N�P��T��>9)G���>�
q������X��.8�;>�M�HdjV�r�z�ےC��25�x
��c�ɽ��a�C�S{M�g��xMBR�p�:�JN@���\���|�|���9VEg�A}�e� L�ȕ��@ڸ�K-7��Ӂ[£����rH��՘���&����3�u��=p��	�s�֏?|>Y�6ߩ�?�/�/�t�`��+�nธZT͡v�c�����6jť�CZyk��r���4?���A�2�O��ח&�6��	���I�7��~����d�����%n�̹�%B���9�n>�طVtxpz�'�h��93�z�2��G����q;��0ă����r�_�6�t�8 ���=��N�OU1����T��Fz2��X����i��ˎ��z�J�_�G�.,��+��T~��\��]�RF� oX�����t3Z~��;to}6}W���	���&H��Dx|P��S.ŉ,�;��G�������֟������*Q��p�6�T�缔��66�BB�NP�	}E�3F��r�
=�OH����d�#�|	���E�qQ��ܣd��:�3����j�E���=�.�E�����٥��#�� �凉�/���?`�����;��M-�-�VaRO�a"vK��r���4<i����="���T'(�G���Y$�+�,-	��:�6Ȕ5�(�����h��E����ƪO��*�m�ZU����Bo":��Z>R�b�Ex�
���̞����(�f�gA΂�ߞr9Д���3��}�q��`$�T�O����4K�2��,��&�`{��$ȋ��ʑ �P�}P�^E����)QY�/�a=�:�:+u��n�9C�Z��<�Ü%�n�q�k/�k�i(Ӧk�f(޽��;ۘ|$I��?���D�g矸o�z>��q����Y#n��,�fK����!/Y�ϑ����3W�G�D�����D��ى�r��C�?�&_�~&36��C-�1f��������{�!�r\=&��:MJ���@J�dݻ0Cm�ћZ�RGL�)u.���M<�о�j��e���;�a�!�U��������G�=���6�;�*� ����=�,nmftC���+��RO#lX�.������f���2[�u��{�a^����+�;�:�q�3;��0/j�F�iG�t�w)\�ƕ?˧u��e�7h�YL��p�	�{XY�v��,c 's��-���h);�?/i�_]B��hM���<8��S ��b�8^�^�'�9�dm
G_��z�Yz"�(�!W&c��jMv/���9��ê�U�/��D����W���f4c+��D|�������}����@�gn8�=����.A�2�JD-o�I@�X`O�$f�(V��
�I��j�֋�Ƨ�'�������	���\5v�W�|�يy��g�8�8?��/Ԏ�h��C����{�>�o~PA�N�	_�2��8�SlmD)����{�^O|��[Q���L�����SZ'N��2��H_�\^���O�H-��ץ{
!���.�-���>�e���&��OJ��;�fn$ ���� E#����9�[�6z��%8�qxw&��7��
�����,�q�ψ�Y{���t�op�t
#��q�O(S$=�j��������q���V���u��mA�Ҟ�#Ov�\��4�H뺲�~������u����M/�ha�I��ӕU#��K˲Bdߌ��3?_*\���`=(&r�F������WX��S�t�ar�%у��Xo�'k^�>�Bfڋ����Ԯ�<}���1���w�jсc/ <��vpώ��6ξ�ʜ 0�(�[}��jO���!�����s퇫U�̊�1c�+��;���Z�o}W��T�Γ--��e�t��8��[�j� Q��1����U�gɞ�??��&�X�W�E�l���X�9X��i]��,,gx-�"|�2��z�����I�{�	�hj����WZ�гf�����"��ړƳᾡ��B���ڑ�ג���z��{�����'��4C�!}��������lØ�^�̴%�,p�����w�<����JU/�V��g-��EG�����UpSA_`+_��@K�0D��[mH >��ҭ�e����Rm6�~w���
���Xa{�Nl7��ZΡ����Vf�6��{)�"u�bxq;�w+��ƅ?IqЮr6HI̲����}�Cào���l�������e��LU�XXz�ׅ�}���y�7a4Gg��ͪhN=�]�$��F����Nj��4U�
�+�����Ŏ-�SE����rh��|�u� 9���9�ܠ�5����u�tX9�X��1�g?e���������O�>�69������W`���F�b�-S� ':����k����x1Y�\�t�K�yS)1�jQ����B��H�k���:A�Se�Y	v�l�V���7��aw���3�)��N���OM;x�p����Ć��*p7I�)�,vC9��������P{�B��>ެ�ܲ
�J�Nl��*�U7��U�u�oqhR8s�\�Z1>��!®�1�vW)w��ψ���zߺU��Dr������{��؍|XаB8��G�'�A]ǯ�+O-<��5Qf��<�vHY1R�����'�-
�NOG�&�pM.Z�$����u5�G�2n����x?ܳ>�Z���, ��}<s4��A�v���˅ˆr�oi����f����.��yU��h�膨�p�S�\��5h@ɩ�<�uo҃���%���M�r�ȷ��\�z绹i���N�ˀ	�仐_�MQ6����g]_��׵�B����aE�ȩRo�T��%E[<��bjyx7"�	�nl(�N&��{v2	�����\�8�%�iđ����݈a;���#j�,�uK�,HEÜluN����"h�ǟ�-�
G�jЛ��j��b��u�����������  hj'�?��3_E�����W(�� ý�-��s̆��9q������^��r<�gy�
S}HQy�E���T^#:�#�5����0�N��p�\�o]X?o��,�1"���7|��X�0����SE�s�F�Z�/����1X������Ou1y؛�x�裑���#�<J�"�1��j� ���5�JO����%+����������E��#���4D�Z.[j2@K�47��g6:�7T�~l^��J����?;�W���Q���"{�1iݱj?���ݦ����W{=����e��):��-ـ>��T�u�L!j&�˴I�9ލk�.�(9G�k��X�g�${s�rzyy����@')ңU���]��m�L+��f�:$�,�k�yT���d6R�S[忬�hX����|U�U��
��O��I��{�Q{��1�Ɍ��=6�빊��\؝������T=���d͎����� ��l����Y�����5iW���z|>~r�[�do��vJ��5�E���p0��Lv�+z�iP{o������Wt,KT퉪��a��6��֙��P~i�(���#���P8���݆a,τ��R���d��7'ʢ�\���լ�T,��Њ Zl뿟<\���Ǎ�R�;�؄8V���CB�W��Vw�N�8u�e��*|��.��G��k�E x�#�A���Uz�g�_�ۓ^:C�h���'f���f��f3ڜ~je�E�����ǟ��AI��+��K��3��]P�3�����d���d��̬��~��R�I܄�m��S_�؛�TV�|�Z ��K�֧�(w[�p9ڔ�Vu����A��g��hH��I�����b��OyT.dR�|��Y�o����|��f��N��&||��aJ=�ٹG���L�9ךU-�ώ�'�SA��� ��ȓC��^s;Ӝ�*�A~�6��*�ţ� 4ˑ�K������O���j���%D8��	����î ab"X1�{��iΆk����ՏK�Ë��uu���ʴ�$I�紋Ȼ���T�.{S����#�5)0�P��:����m�kY�����;|���"�r�s^Ґ1��r��_���a�����H����?��Qnk�]���<9�7ݐ�0��xA�Q�iI.i�,�\#@p������ݎZ��߳ܮS��>�Q���9�d�p���m0 ��o��齥��G+���Q�w	�!(SY0�j$���}��h4,<�U�)���k�Yy�*V����]lI����)h�}��u��{�!�5OG`�����q~�4ص����6����|�P��p����;2(�����1M:hJVCE�UՌu���zzl����zS_��%�4X��{���D���C�<%agF]<9�FFaE/�;��ԻgǊ5�,��� ���R���ۙ
~����y��g����o��d�%>�B�[����v�W�w1����NG�
X�[@l��el�sdo>9g�{�W���\�� w�7װ�M��.ه}C�W�j��-4���l���Ǿ�~�P�y�K�¿�}��O�?�%���BK��.t6[�}C4dk>*�ౌ=���5'ڛ�'�3�o_�Yw�i*'Y�O��v�q�
6�&X�!D�v�2�z������>W�
H]h�e=ح*�����y@o�*W=��M�Y.g�Ԭn�oҵKn��!h��F��|�Ӂ�8�+xk���'���4��P>խh��/qN�O��s�����cto�� M���l����h@v$�=�NGa
7�,���I�-W�BΤ�TJ���w�B��� !�����I��x%87v0ȅ�fK�|��5���)q���#kP��e؞��'.\�	�H�N���m�N���oWP�~�F$�M��gD����誣����(* ��#%��H
�����t) )-=0��%�9C��)]�1��90��������:w���9�sat�~~������a$!LB�e�(���2��;Og_�5يI�x�r��p��w�]�#&8o���肆��U����ʼ����gָ��}�oe���l��Y��U������G��zi"���Wh�R��`�2T���ҭ�QB��v����jl�m?�?��AW�G�;֏��F�ڛ6�*�1���oZ�u?�eTT!}=��ȩ�-�_NT2D�b�z����	w�Bъ��Џ�������������nm\�x�G8��T��\L�e�ș�U�������zٜ�,yd�".1�=�����.�#��{>v�����ߟ������ME���>=�����������׶��	��ט��ݦ��"[�vZ����8I�ra�h����G>�ϬN��w��T,rMޞ�ӆ��YOJ4 V��#ⵅ��cE�j���YD.�w!�oE5��'�3G����gŮ���ؕ��t�RYi6���R���PE��X9�I7��z��s���1%bR܍�;���^O���W9Dqr<�������ۢa�I���>E|�[����
L`���l�*����_>_�֟������F�W�N��\㗞CN��B���/�v-���1\�)9d� 2ri��^WعM=q�	�{F�D\�������jo�8/�ɫ�^{��V�l�R�M9<׀��e�s��p־bƯ�4�KTOl�5�"9�\�������Q�\���j�T�l��G����9��N�_��n?���Ӽ��!�,1d�0��,�h��X��m�ϨG���&��Mɜ��������@�2���m�[��I�7��?�PR��J��sG;gT�����א�ɍ�k�W��:e������g��*�q�$~�
P�ؕb��o�.�&>L�?�\�?���JmL���y��*8|r8��X՛�����Ȍd o�v���!�ωS��ヒ���?.b�}im��7�g�(5�ܯ��
�O���;>���������=D��P^�5�Kl�V]q�˟�7Ry p��s�tP�iSE턣Q[����4�.�Hs��TkR3/�XJ]:�וu;����Tq�;op�����N�i���j�!"˖s�:�4 [�W�,,2����B�B�<�FR|�\=,Y~�ז�6Qc�v����A\Y��]�;BR�0����t��-�7�C�T��dk�Eȫ����¤�Nа��i�s���e�L�㪞���[�\�Nn�j�]���̨ڸ��+i^�FM~O�V�!��۳��`���+����i�"�f�oj�;�1j��Q9lg����⺤<�_���
*��s���s�2��)nWɒ���1odȰ*8Ь��7C�`~��H��\��D����@��4X�����t��}_�['���	�5��k��jj�V[�и\O|��ڸ���@��،���Ϋ�%0bB1�k���^�׀������1��ڭ'���=��9�6f� �T��;8��Y3��ع����U:Q�X�v����0TA
��W-J����\a�fr�Q?0����z؉�8h�+�I�y���;���QV�k����������:�B\Xh��Ь�}
����юv�1��`�`/���W;���hy�)?�'�I-�y�}��R�D7q&5��`֜@�j��-�V�n(���d?S�,8�7%F*�f`��H�������f�M�Y{���;���M�+I�hz�85ã_��>�+�r��y���3Oԋ�l�x����*4E�y��&|w���<����) W�X[�I��2ɔN�����q@;t刯��3���5���u���:�;��u!k�ʺ��P�7�rA���!�4�KWJd�ǌ2=n��"W��~���ǻ:M�F�{�%��6X��(�z�������}bRa�hp;��T�,�8J@͂,*�6�>��hC�ǲ|��G'���d������e�M��;���[�"J(&�3]syW�آd.|?[��_r��F�}���~'��!�t��jp8V��w�KV:����) ����V�4�|��UBB�^��e5��%��>���9?&8~&Vt��ƏU�{2r�����sJ��+���C��,���G�۩z-�~�8#}����,ܧ>�L1��ꘈ�Y�����In+,�[�s2iv0�����"�EN7م������7�5֚�C#j�06l+���e�<oFx��Φ*������m��*��"wbSrYG}΁�9l8'��Q��7�ׁ4�(�JW��_�X�E�������S�֤���J[�����vo�XV���>�5�U�d%(�N�吙�?p��~)���zq�O'p�H#+y��dlr�Zl	��Ҍ�#b�D��$����h��W��`���8��s ǿ]m#�Х,��3�Xm�|�����~`d�M_�Vf��x�>��;[������_�S,}��=5�� EA"���67v,D�[�\���	Q�S�c�Yk4�!-r�ثaͫk@��^/͊�tO����n��u�o(�mp�j�mn tP���¸� �:X��o���0��6Q���w�w��%]Y����5 (]q��Y%����DǦ�hƮ�doo���4��j�l�i�i�zb�w|�bޕ1�9��̛z�=����9��`��[�l��2�y��ک��_�]�t�An�X��g�P|$�-����y��M\/̲.&�R�:��y���lc�~�a �k�Tv�ߑ���¥�,�/��_�
����a�|�'�O�$@�����p�
�%�̤g!/��'#蹈i{�:���T.s�83ϰϜB4���9��ʵ���Z3I��������q�����)���Pgm\G}%������A�f�j��@�`?�-ת�i�����Ħ���y:=MT�N�@y%�>�Mq+���L��,�#n ����V�J��l�":5�ц\3j �WR��-;�1W
O�A_xfB臆��ܗ9�Qw%���~�%�.g&�,X��D�CmF�����4� ��8_���@��x�/,K#�O�1F���	"��Z�^W/���6��L��?LP(w_^
�y�uu���b��o��X���乃N��@�p���*��Z|o�@����} ɥ�'a��+C>
�g�����v�/�Gz.
����A�rA�?�7�}�pI�d"�e�oe��U�?� �a8j�`��c��p�bF�PS�F��ٮ#�`���[A�z_��F���������{��B>��q7���e����O�(M:'=��i��6�I3���V�!��z���o�<Y�wN�ƽꑣa-f�+&݉N�?:N�����3�upT0!�Ś���]�x�B��?�B�����We[i\���嶙Xx�G�*a=5���,"��s5ӿ�q*�+2����Q.�����q�I3�o��-&��̘<��A��qMx�yF Oq�#���^�7��}챪�]�����8�M�ݍ<��Z{����'Ȼy�qd: Y|W�L`8�i-��]�z͚{V4�E�UL/� �e)��GR2���1t����ƝĪ���Q���u)3%�/�$�*��:�a�
�bI�!��Q�?���
}��*�͍w�_otoΒ{��N���l�!6�@��j�$���R,ak.�ɠG|���u���-K�E!�9����0::�BD<���1�,�1O�m��(N�Uǆ3�~��ٗV!�uw.��,Vie����ד:�7#_%�7�����=_���ʵ��8���TՒT�d�~XK�d珍�����'1��ĩM2ͫ0m��r��3�U<}c�n�$D1Z�\�I�%�H��s�p`N�I&����t����X��<f�B��Z�$Fᗖ�*u��F��S�R�q�:�Ӹ��� �Ͼ%�l�lay���u�f��D���犒����Sg��W(�M��dK�%��~�{��?]n�%���8/���@I�F�ƫ�'tg��/2���C�_@k��-l�1H�m��]%��{��P0&��2�|��؅����y>���B����VJ~�������|��e�J�颛t5�b����U�*��X����2�Q�r�(w�/MI�s@�"v.��G���;UoM�
������_��Xْ�)�q���e.)�&B�]����܅^��&�+8���;fv{%C���A�ȟ�-e�gy�_�1����_�W�ōjmA�`�}N!ۙ���&?�?����E��Tϊ�
�Y�UMBd��Z#�W�
ԉCj�T�.�>���
W���\C�,Y	ϳB5�ԍ�SƁ�wO_9�t���{��T)��

��Mo^�P3)JgN���H�{��fJ�I������V?�%�am��$��U�H�jT3���_{%�9�-�03��U��6s�5����7AL��*tg-�'���`���g��/O>��A����q��>z��Jr�<�4onؐ�Q�c�]�-Х.�7b�N�����f�ğ^��iYd�e��(��qɥ��vY*M��1��4�
��߈��݂��W��dD?�w.yc�[ЖڔB���؏l]=�'�9���ժ�|�WzH2�����E�(+p'�f8��h8rй,�პ���{V�nz�������R����EQ�գV��������1Y�?jԋ�ҵK��8t���w�Yh|��H���8�@_�~Q�e�{:�Qh��ZQ�5�an��ͽ��MC� �/.Zm��K�R���;}M�ه�k؏f�<�Lo��S2����fq3��T��>�>�k�B�#����5�`�߫N��1���,ޥ왍:u�Ya�|�>(Uj ��؉ݰ��j�{��'�;�$�����ߠ�ej��H�x�I� ��R�`�3���3�Z����i'��:g���_�k�Wl�����-��)	�E��
�	λ���f#J$��4�\�P;�@6Y�U�
���':d�j��� �P����LJxz�p��C��7U%٤���P�UWOm�w%̹f'���o��}D�����[H�V���h�083��.Φ_3v��?*۔_wi�R���z���p���f4^���u�5��XE��s�ȯ�w����y��b��� �:�kLuZ�%��p3��u�����#j�_6lGok[k}m�b��vv�����W���D�pʙ��d�tP�b��va:#[wrgřj��>�j�wc�x���3���ӄ|)m��՞��Q���<�0m����#b�4�v��.��P�O�2LJG=�h��&z}��H1�Iv�e7Y�{�ѭ�8xu �����O����3�0\e�~+z����\<Y�sR�Be��S��O�0��.�D��z�������c`�s�}f�bL�	��k'چ���z�m�Ȣ��C�s���2���5hx�fxP���p𤱍�
S6�]����'�Յ���_J�cNd�7��Ml������R�T�	Z�p%z�ͦm���;`s�sC��E����M���6E�Yuk�AA���qb�>���f��p�>U���h�3-�k�Xm�&�w%�j�7���ٓ�:�>	j{�fy?#�^���}. #��Х�����Q�����^eu;�W}��<�Z�Оo/�}G��$���=���J��zX���0��P;1�=}��
�2�$v�y���r��׀OѾ�x�E���彅���xEw�6�"9�%��ҝ��7���v;M)��G%�X-9m�܆�hCi�h���X��#�����9���ȯ���|FF���O����^����f�!�2�&���p��]PZ�k���d�<�	3��/&e�E��ы���������I%(�p�ƿ,~��\:+�O�?'&�N������s�����J��]��d"�ijF������~YXk���M�DC�f�O$�k��Wkk�n%�H���*�-:�$'�p��s����3�D���Гy���O6%Ro���� ;�Hk�o�5��#�>/7-t�{�d+32��_�G� Y��`�>Wm�"��	NJ[��*4H�`Q��f-k������YS:`��+��e�i;ܙ�T��
��˾�E�L��,��@ 3�LP���`<���N�[�V��l�=H�ٛo���Lf�9%~B����y��m@�mV��!��˴�l"&b�c��(��*e8hu4� ��(�ng
L���<M�a�eWP.�8��cʗ��-ZA��;u������_Z���NC�\Vs�ne�[��a�έS��h`E�����^Ձ$�˰��g����������fs�����6��
��m���*G�i�M�w��J��3.�}�<�b��@��X���2�FP���S���U�����R��o�G���ςn�:��k����=���Y�׹ۥ�zKC��,���]O<> K����͙�/��(0�k�]��/lS�{��U8C�9��3�V��<%=��c�Toi��-��p�?���!;Cͨ�$&�� �.	�m��:��+���ȑ�{;.w�t����z��E��P��E~������Oy���o��l><��t!���8b��':>
D�\�_J{vS�v���\u�<����A���עܚ ��[��?�t~��_]�ԢW
�)��KW��o���X !?nN�ؒ��������LQ�s�/gij�w6o�V��g��{U�"���EAۥ+�K��<���˼����v���mq!a���7{B�W���%�#�¬�]�a�m��j�.��y��M�o!jS<��rt�Φ��ى����s�ewl��������W�6�9���V@���$:�%h���[��2���Hxba����A�IOa\�q��ߛS�[�ue�$
�hLpG��zs��3|bq���?:/�ϫP�S)���^r���!n�r�A��,�ߘ�Up`iѥ��"��ybp�i��%�l�1�V�s̬���</6��F�c̺h0�Z���%?��9�s���1d#�q�(*�K�����I�)������@Z+�5̒�(Z�U%s�i��P��T��V���Pkx���P��B�����姈S���rZD1���*7Og�ьk>7�������)��:��5'VʕW���2h#�G&�S~���~��%��o��+��m�X��~I��������we�]U?K�=���92�nm����ms@�l:\=_e@a�Y�
�|v@�%%�lGJV& Cq������{�
O�-�[�_�vVz�[���N���3�1���m+&�M3aK��6L�k�8@*p��;R>��jGH{��������¸^st��h�N���8ɟ�<��q��c�j�/ٹH��Yh~T�X���%���0�hʜ�xlj��Ƒؓ�4߻%7[R�|�F�5��R�)[�y2sr�����-H��ā�MaXX�
�ݾc��,�������{ �b�v���]l;��y�;����#O��v��|������Fkr	�sL�aԊ5�
�Mq"U7S����R@5M��T�H��;��I�W�u��{�ޕ��י����7W�������_���K�l;f��nm��a$� J-q��A��l�"�(q�������VS}T��t;��/�~������s�!�Z���h�ֿ��Ò���"�g�A3-mv���Z�ϸ9���i��SV�e�hw��Dbx�%c���*�<%t�c�/'��8�@���f�:�R�lˏ�W0*�.�ءc0'b���	��L2`�k�iq��V��0$��p���nhPu��@Y�}�h��nWJ,�.��?��m��k@~7N�.���;b{qZBU�+:�z�v̇p�&��}�^ڬ��L$g��q+�������~=H����"?�"�~��x��W�&a%C��Č<c,(ߓv�F��h�4�q=� .�ׂ�ޤw�܆�
nG6��	'ro@�/b%���pX�[*f��������F�QobG�Y�_]����X!+ts�'/����o2�����1X�LV��k��Z�Ϲ\)����{=���b+O�FN�}���
NqF��"�~L"Rұ���H����{�
Y�2�C~�3
��\���!�g\�
�2�Go�w���g!����$Ӥu�z��ֽ��j�?�[�5 �H�%n H�G��9v9��uq;[��,EJ�������q�g(��m�i瓍vD�d�w|m���)D���5@�kc0���{|�NV��'�&�Ŗ�!��������e��|mg�Բ���#��-��=����˲|7�bm$���
�����.e9��twQ~�6e?,e�m�i��1�k�G���!�{&��-l�z����.�D]��9��6�4J4Lf�}Q�G@���&��k@�&�fP�ͷ�-�f�Q��}��z���,�nkNku��^��h�(s ڧ0}q7W2�n�������Z��g���3�	���4	3e�!���傟'7N�>���l�>;���x����Q��t�d	-�lRsU�[�VX��O��e:@u�N�2x@�WZ��+��҃��9Q�����ڥ�t
֢"���Јp����kcZ2ZT/V�(:���|5yZJ��y �����V������:�Z�e�g.��[1��c�]�FYL
^��_��e���Â���nu�|�GB�.��ف�J�7]/�e�[kV�+�;��Н����ą�c��=G��=�H����+�Y��w?x�)�߇�h_���^�#J�x)&�����}nd���������
�>L��݄�5������=����:�%�>N5����=�I<Y�U��5��}�M���h�0*��9`#��d\9˓����+}�;=t�� >��l��GF��WWtVfw��,P_E���ԟ�5�"��h6R��PN��E��G�/0���~�@k!�A���/��Oα���h��%�\QA)���B�����?Pa���C��y�*�?^[����)��y*l�����S��+�;mt(�,b%Q�����uk\s��°׻�.�B��s2b�=v8�SPkT�2���sT8-]�rp�M{9E�k���������{RV�eZ�<r�~ ^���U�Yr�y�/+E����Kֆ
<��j�~D�bn�Bո��������=+ݢ/*X���8��.��(�Rハ{��׷�J�p���NB�L �*殡J�i!E�L�{j�+��E鬕$!����]�̯O�{:�K��nٵ����j9G�n�WS��[Nd���r#L�)��?��+����枖n�&z�F�[��J\��V���@�E�*}��{|��q�p�w����,Lf�s��5R��v�>��d��3��L�tㅴY�?�$���셴j����Ex��".�`�WRX��'d�]�^��?�'ڔ��>�����9ϻz,�P&>���\tF�[U5�}r����39r�6|�er5�R�^�3��]�ݼ������薣a7"���m��K!�O}|CM� z�r�>�[��D-�G�JaD��)���v�;��ȍ����T�0M�8"4�������r*[��N.�q\�_j�Qr�.�������n����\�h2�vͿ.��{��Bxd<������"qiBu�-!����l��~?��.�n���v(-@���M�tW�7�����(Jx-��x�k@`¼<Í7 ��LA	��o�@�jv�D�BÇ���ΰ���L�r�?�Yk |q�CR�F�b�P�kI)�5��P*p=\1�ЄXc�k�w����A��s5bTo%%v��XM��˘TE�D�7���=��˖�-�����f�+|�jo��z���A���,y�)�=�=-�W�0}2���*gȗ�ۄ#2x�H�C�i�� ���0@����r�������ܬ����W�����ZXO�ܻ\9Q���T�+���t+'`�!��.y�Y�Oڶ�[Φ�1w�2�I3*�gkGw����r�f�b�5�9���Jd4i�N8ֿhPZ
���U��:��(סa�T'ܕѥ&CݚV�$(��c$����K��֔����&�u�wKCc!��vL��d�W�2��8���Ծ�g#�ăo�Ē�?�,��8�h���D^��q���|�Ѽ���n>]it��X��Z<�e|�(sL�?�j�������Hϧ߄^Q������"N�Z^��_�V�HJ &��-F�����ܾ��E	��c�m/��[�H^��蛡ޘ|�KGP!j ��7���R��f����o��2�p�k�R:`.2�"�e��v���q��T� b�{���s҆/���ɴ�v�����o-t޾����tQ���A �qCs�Q=(�T��"�@g���b��]��t�\��2�N�>�����Tb+-��!�=������/��-�Ë��T�ȟr7r��<����%Y'4�@�:��2bzu��^�"�Oq���V��6�Iݙ�2t�(A����1�S�7�W��jwU�=	��E���&������{���D�@�߭�>]�$:����lz@�x�@绯뇉�9i`�Z�V�]G>�r�.Ѡ-���~bζ�r�]eV��M.�+?	��"��P[09�i.�[f���]�猑d��9T�v�<��~�X�x"w��D&s�<4�V+��?S�|/��Q�}��^�/gF�eK��	�w�LuiZ�Ŭ�CB,�0�_<Z�'��ۙ2�s���T���~@2@:���Z�Ж�̚�����(��}y�a�ƙ�"�ۣ楡J�-틊��hl�[�3a.�����{c��ݻh�C�0wk�c8}׳%��[�>n�zT�m���su���`el�ȹ��u���T��B��DUg��Y����T��RF��������)���%UNk��x�.�Rx���@	Z�S�qdA�,�m�q�Z���	�!3E����&U�(�c���ݮ겂�Qw�c	!g���m����T�B[��J��-b�0��IȻ���ڟbӽ!�g����O���>�S�u[#�ȉB������q��#����K���矃���x��:��"�8r}t�y�.ŉ@S�.�u��NVL���~�AO>}uz���q��Fic�QqNg5d�z�i?Tf������}�J���^��GšF��tI��T���g��Ɇʍ{�lb%���2�� -�t�
w[l��^с��o�t�ݖ���M!yW�����X]�=Q�!�ͱj��p�꧋�\$����)����_��ԓ�Q
s����^�s��O��w*��se(�:�f��>��$�O>�<�G�� �}�/8����X�E��Yg�͛C��7&�[c$�Q�*إ|�b������*W���q�����*����k�m�jz9��&�,4TA�g����T��'���!���"Z	�����-���.��sb��<q��Y��	ی���}��f�O�����]Pb�[���t߰.�l�'��|�B5ߛ�.��m)}/�[&[��`ܺ��bKF��&��kC���d�4��V�*��������D�&�y�
�F>L���
�HH�	��[�ѐyM�2�<�Pu�5����[B�2p�rl �mF+s5����a��}$�\0��6�fn.�E���6�C�R����z%���f�a@5~�\o��i��kJbVY�a�C�6�f���$�iN�m>w��0,��QC5Z��:�A����a���˭��,����5���oN8g�RH�d~��������U�����R�*�c^֬�h�t	t�i�]M�`�ฮ�G�	�L�G���#(�����_Q���g@����d�.��sZ?��}r�U�B��;��AF&�g��������T�WV��Z�Q̙N�2�q�Z��5�	�޳�yk�@��UtM�$���M|�	��0b!�6�ELHe2���#���"�2T^��E���T�����$��_@���F=��&�%�v?�s|Nb�П<c9�I�
g�Y'�$j[�.J�<���;��a�����0�b`����9����3��5��k�_D�MT,j8��x?Pia�է���C��!~�-��XD)@�e���\3�χ����F�)/�3�Fxϲ
���B\���f�b�8Y�YwYAo�lӍ�\�JP/mD>��>���ŗ�,���K�59L�U���e���!N�}{l���3j0k�7�dr���yXV���4�ڂ�,#z8�g�mr���k���(��gV9��y��?�[�q�i��xH����q��tɵ;~��d�L��i���Ԙ���A�
�f�l(��ȜB��23����0h�1lA�X׭�y���܂b�EA��U�k��=>�D%����LvgP��!����r-+T��m��k�?u�IH�I�����.*�d�
翿/4w�
M�n��zQ�%A7�D~_3��1��0a��,�>�>�)(��s
��<"�)�{�]�[�]�`�(srm��<��Mqy��3��Kb�L�MSv���׀z����[�}����6��_*�X���:��<�\Z��Rn|�� K��;A�[y4һ �p{A�"v9+K��oܯ�3�i����B�1.1f��fWڢid�tB�
LY�?x!|�'7��'�"�c������{zo���F5H	!e�_1��l�hҍ��zt,�8�ÿ�2ҝ��5zס�C��4�s8����=�/}ǟ.g�r ���d�b�fO���](D׏�Q�#i�yɾ�w��׀5�<��?��0a��{Is�dO����-�)������RA���{�d��K���NP�}/���O�C�z������ޖ�N������ڠ�-�1�:�.�t*7����28� �)��sgg�>U�eK��yT<�~�T�������W�=5O��w�p���P�}��Ųӱ�^#�{����I�j����ퟻ��R;��,������6�U?ГWNw�ƌ��Q��ȭ}M���g�.|�j,���&�p߻��q�;(��?߶���f�vӶ�焼�j�t\���y���ӸkDtJ�4X�G�|�DcU��=�C��䚮�����5�#-����j��ӧ�h����兝k ��$ ^��f�]����Z��������3������diz]R�Hkՠ+�?P�qv���c�}�ĺ{�zvƤ�������"�6 F4K<6�ş�����&�����r8�V�(�΃�U\B�z��x��>~}��g�z!d��J�.e�n�U���Xk�~^��ʄvʃ,�����h�{d˛Uk�	='_����C��N$���f:?����]�
;��̰�J��xq׬j(ya��jw~4jy�j�#&��r��v^��:�{eN�����B��yN�l7����*'4;� ?�HM�Oo���(R.�7��0b�%X�۞�	�]���	��a��姦�z�p�Lr����?aƥ����a��"�1�{�۫ 2h(��m
M�ח��z�B���$���d5G����<Z?T�
q%�9=E:�'�z�I��d�fU��z"���� �� K�V�'��Aj�2�1J���F��E��p켻�"��W�W�%��b5�Ax�+B��R�{#K�*����c`Tʧ��٤7��o��y�#u4���'Gv)��%��cw�E�x�w���>-Q�dx^��OTo<kA�Ꞡ���ߘ�}3�t��&�{�-�\D��G�#�5�L��KLL��J�Y��@{�y�&����]ѓ�/�+��߰&j&�A/�݉w�Q�KC��av
/���Z�n�boMz�RyKV���G#�+[�ןU�sJj�M/�e��&�6�:拨�Np�=sG�H���D{+��U��([PD�O����ߘ��N������H?Uᤈc�NU�m���u�	�nLS]4&���1�9���hs�k��$�{����U����Uy��S�&?�{e�^����ʾV��Y���9��AR����.T���J�I�+֚�E��8����G��q2PA�����j���� r��[t޿���o��"�a��η#�&(��D�����C��ֽZ�hP`�!pԷ>Z�UCݩ$���Y�'P��8Q� �J���į
�ě���"�m�V<*���_Is�FXUv������?�����_\rƛX8"jAY,���{�j����1$T�'�ыSm��(��z�����q�����/�^�踎?|�{�	U=ly1�<��љ�#���&+τ`���Jh��?���І���\�y	J�m�]����F�~�PB��I����*!<�l��E�}��ю��P�SYε�a�5_qb[��{�ݨ�)� ◽��:纃�<�ӻPi(��Dȗf�)%�2��M���~F�X��F���8�b˿fM��w�C��4�+q����i���P���W�(�n�噡t��f���y��+c ��˲�&
�f�'Ʃ��(	t��'`�l$���}(�n;��(�1���~5��0<Ѫ�w�i�0z��X�ء����`T®�_5�J$�SW݋��߽>�
?m_,9������R��Wb��ѱ]j/�^�(>=�KV�r43K��,MX%� ʗ�炘�|���x݉J��->�n����qa� ���F����Q��P�6/���ш�Wh��m�_���L��\M�`����@�b�`�#c|��u�����q��I��gr+�C���A��x����1T�z�==&i���:k�6s��v�xj>y�Y*Ma\�u�j��������R1 :�0OC��H5�i��;��tǸI�\�ou� ��ƾ/X='�����-�:j��p�1�u*�����]��'�OM~Nx�RE7�v����)VZ��Ԡ�Б�������e3�D'ᲊ�o��N��ɢ�/翅�Ŧ�8�L5��*9��

�Vp���}��<�2"��{���=f��feq���u�"���M���*��u�'��[��\z�]�w={Γ�*V�-���`�?7�y�=�֖K�Z�K�h�o�؍2?�0e���W���z���}2���3�R��x�s�+k��jH������Q��sު~5��:?���r���KP㮖��W]�����p����j9�m�����M�8X�)c���d$J�-W��S������W��K�Eb[T�	=ϴ���2������
��Mx��s��dEpq�S��9�~W��K62�z� 2}w��ڕl�����kd��<�t+���L7�F�	pJ_a3�1v°J�J2�;��Xֿ���{�(��U2a��	�:6^j��Aq9�����	}���:�\�q67�'ݟՎ��X���8�M�%sv���8�C������&���im�'�܂�-iD�,�-��a�?|�O]��XǛ�P�
}��U/��`#�­|,6�O܄Zԟ���v͵�����XĈ9�8�YÕ���a&vg�x�?�,��J���ٌ+1��E|��΂��%��w������B5c[���3��Q*a�jHUܨ��°���l�k@�'/?�a/�������P�X1W8S�)e#@�؞���G����rϞ�% C��0�G��:1o�O��eryL���c3M����wB?�Ǐ}�?�&�Ģ ���}�J�?b߫,�����*$\PF�(h����y��u��G��poG��)���i�
o��33�2�O���=��#�q{D��U�G���}  �^�h��Eo�Z8�ۮ~�'�o#F�=Y�l2�r��q��fN���,hM)�EH\�-��g
��%�����8�R�ݕ5�
�'�ĭAS�S0R�b�C��>/�\�x7I_r�3`0���ïXĎ��r��"�]��� gb�� �Nc���5 &�}ү�e{d�}@��~��sZ�IK��ExW*B)�U�m�,afP#'XEK+�À{� B�^s�9�o�-ݱ�Tw�n���/z����G�*�����?����Ewk�o�D�* �C��M��(�ˇ���S��F�T2�~��*`�;%�Nُ;�i��Y��a�U��1|,�*˨�l���u;��`�	Rcw�]�,ŭ��	|��� ����(S�2��@	m�Y��Y�<�k��	��
9.�=�5�)Sj�ָ�v�5�U���t'�$n\$>���=Z��Yʁb$��!��.@�w)h�k;@�W�d�HP��Y�W*���:.v�i�ͪ׾Y8OQn�������6ͲnS0ގQ���[^M?���i�| Lr��sUU4��A�пn
���ɌMk���^��ob�uLv��rY��5ط}�?�b��*��#���uG�����*m�*��-J͖�#m}�h���� D��HQ�V�V͔�+��7��BbDH��������\��>�g��>ϕ/�i���sXV��h�B�Bt��X�_����r�Ұ�}�Tn����|@&�,E����T6���ϻV�c5��j�w��S/K����J-�ep�1�C�0Aɋ.f�p�b-�+��f�*�B�GU�{�l�8�|ܜi�x-{�=�L�������ӳ����=!���rWɫ,y��ȩ��nL��1B����a)>9&p[����9�8�'۩:E+�	g/��&(�%�r������6/��yj����<xSI������M�Lz��ݢ	�F�tX����'��;w\=:�h�Zx�b�/�.��<йǘ���-����kac���G�ώ�o�ɿm}������,�6�ݼj�d��ǒz���ܤ�/z/\�]�o_��|G�"�c]�7|�%�u��dL��֤�����C�]�����J��(����$���>k׺����%�Ŋ��Y�.�߮|�6�&OW�@�}l�I�e�΂E�#1�	��D���Ŝ9 ���4�5�����B�~o�����^��u��bR�^s� _H�<-"�4����[��7::�{Ų���k��߮|֏B�JDl��Y;�h�������b�e�>?�����ه,d�dѶL/9|k�l�p]&�=ڳ�U^n�W2B�W�Ԋ-,��V2�ZTQ�c#mgB�����ȃ��m��'�U
��K������S9~�'��}�*��y��o��Mg���qů#-C0z�H=���ڙ��i�-�4�|\���+2���
��@%���z�y�n�Y�By��|�X��:�����}rT�pW�DA����X��}��S-�S2T��Q�>y����1j����ac�	�j���kٟ����(S�E6��A�o�.쮫^�CQv�E4p�dӯɫt�D����R�V�b<V�f�4��oݛ�q�!����g3�L����6������*:%"�4��F�6��9�1����[�F�'^�E�/F�#��2��BJ����
g6*%mX?
�+���<Vx��W���L|���Le�{s7�|�L#�R��Otg�\���*;�k 3A�P�.��p��q�0e���`w�&xGc�+�����n򴻭��Z�s������T�:��D�s=,rc
�5��H�mb(s��U&0���F��p�dh����ݒM���@9�4�94�����tg� ���e�)Պ�"%��M_ğQ2������{�ag��R
UU 6�5Q_HSM�W��m����Sn>��r��"-뺮��-b�h?�A�j{����<�i3n��fvm�7�$���F���ӿ����;�y�v޳ܤp�?�X�),�19F�\�����/����T�N�󉧷�1�j�������T����+~yL���jL ��O'_�Ltl���<Ύ�lw�[�����[_�; xםp57�p���O�Vk���w	��"��M�{��-�>�9DT^)��+�D�0)�����H���%�Z���]��)��`o�r+y��!ZD
ߎ���k�H�p x���a�CvXf�] "]�O�<�Wj�x���q�yI�c�˫�q/�d!DY�ZYz/���%�F'�z���dH��i��5%q�(��g����w�2�.��Ev@S��	�|�Ms��J�<�����q�Q��[M�9�D�9
:�Ad�&f�w�c���eLB�ӟ��E�y�T��
O�ȿ|�vYszG�y�>5O�~r/M�@D�؛�8+j(��Z��o�o��0D�~��h��g`��f��(p����-�5�zp]�D�������W�Y��؉l�ۀ�N����1�J~tL��n��j��fI��\/S�^%�?q��h���Dq� ��_8Қ�䋞��=۠��㢜s��6CP��bk��Q�j׽�=���RgӌD&g�E����&�]s���ֿ��S�%����#��]���� �t6�(nw e��P>5f�s.�z����*�kz����B�1�Dx$('Q`������r��kG�p=Q\{Y��Y�G�V�M�5&�P��j���">�S��T{�z�h����X�����H,���?�4�`�_?�m6{��	�2\t���N'�oM���)Ȥ1m��}B�B�H]���3��J��`��[v�x�����</HE}btf\��k����#�2�'���Y[����BaQ��j2<M6���NYIZ��%���&*���R�����:YI�2AW@���)�j�\�2���&��~����y�������T"*D�(�7?���h:�S����im�l�r����$�UE��ȴ�=Ooo�1^|4z8ҹv��C�]�DD0a1-PN���EyJ��|��f[^�����L��c�"����nn>?�V��H�`��糺L��CW�A�=<�|���D80)�L��P�ӎEI��o�q� ���Hȏ|+b�nR��9���X7ν�+m���U�R�*�c�!N��6�#�μ���5{��-���~ �����*�ω�4���Ğ ��YE���E����{w��#��eӡ�m���׉��0Ԥ�h��P�$�*Q��5�J���qp�[�LFtN�07��a�`����q����5�'�hۄ� i"��*2Lp����>������0��xO��Nz�#��|�����������8�瑕U�Wf{�7[��h�dx�숬<���׫ޏ]�+����İ7T�'�s� )�,���U���t✔XR��υ����0n��Ǌ�ֿq��b��Q����rb(������go'U�]�&i>M;�6٬�B�.w>�U�a���1<|�z�Cڭ�x?�j|���t�Ȋ>�_b+H4�z�ٶĲ%aW6�"���g��c�H�u���M��������G��"Ä^�[[mړ��E���,�k�����d�����[鿡�n�+�ƃR]|�xbG9T�#7�09�q�?��0��D�B@ڵ����g��s�!C�͂	��wٰ�6��6���sD?�9���R�ؒE��"�x@{����ߑ��۞EX�������}���_������ٳH��;RF'ϙ��!P[�'��8�'�}k�C��YȖ�y�iE#�q�֝��$@��육����6�a;n(�5���.���2Ƈ�C�;|���#Ē�hB�v6�C�9z"��X�B�j���.ǂ����+O�ƻ�=p�av��m<��$z<�>払��=[�`��ؕ�=v��!��GV0m��c�3��H��N�IT���	���ӈ�p�>��qz �I�W!���^�"3بC��L�;ᵎ�1 �B���m�a�"+�]��$�O�q�J���9�a������G~�A�_Q_��hV7{ߑ�b�ʥ��M����/��<�l.,��ð4����Ei��t���~ຫ줍����:��-�N3���Hz�w��S�����w1#��D}��'��o�-��-����L�I0Wr��|�M�o��闔��n"����b�K���@���Z6���h,j�!~��x��P�q��4���#c�PF]*�p����졑ʫV��<W�~�����A�&C�@8�7�ȸ�/Hpl��ɤm��Y���?�w��Z���@$�ћ����^FYW��sx�4�
�w,�SQS�CI�?(H�"Zq�t@��{Ff|�h�N�V՛��Kc�/�oZ�P ���.����<l�ޏ+%� Tx�Ds��wݏ���w`z����#�6¾�2tQ�@�/3Ck�E!��j3o��0�s"�P�'������������u�=�u����ȵ�
�<�6��X�m��[�$3$��:�����a�EF�,/*���Ю�l��\����L��Œ�٠�lϾ8��0����ˁ���*���ܔ��S��˽ݢ���
�+����U�q��}�P����YO�@����x��ϱn����� I
� u�
`� ��XN@R6= *Ax���%:v�o)s��f��md�`n��99����)��Wv0��� Z]V�{cC�#*{��io>Ucx<t�[���/$'�������kqvf���t�ߠ�c�ڊ!�/���`��������-��?i+v{��TQ!���������"Bk�J�I���耙�ã���{��?U�ހ.u� ���Fvg?�?0˩nV�`���S
��2��-�$�\4i��%�y�\�6�:~�[R��>���N�P�uƮ�YI���a�6Do~Q /"A���%K��mZo�H���S�}�Y4��L!�ы�Z.#4u��S�����ha,���ʲax�N�!��y�7�d.�!%(�.7V�����׊ڄ�F���X��x��2�/)ƨ���x��VYX~��A�#h���}T�0���_�ț�����F��~R-��|8a�}{�a�k�E�+���g]�����K�^p!��j2X�8ڦ�8�I�#qUlk��Wi>~�\�u�tB��j �xr�x���Jxl[f����}�p�+��s��g�zZ����UQ�bL�mR2?�ycM���/����|A��5�5 %�r��M���4�m����E.y�CJEm��m��2��oB��ݡ]��Ë��%�_���$O�Gvk`�Rm��M���Q��
&z���ō;_�!N�q��C���:�^ь��*22���t�㛵r}"$?�hw���6ܼ�_C��w�|�O-�{�uAY�޼��g���T�<��N�Vvf�F���.�v�@S`u�f�Ŵ�]��b�b(r2�Z2x	��X;�9��)Oo-�;6���G�e�v�v:�J����_�}��m0�i�ꇧݠ�mh��f���iA����E�(Ah�~Z���z���Q��tU`d�n%�&�� ����)��ETZ�i%;�|���	�,Y%l����c<�}���:HD��qI���K&eIpYl��?�] P�����/̿����p�o�YX�Xjr(�`O����_���%�d8՚*��0��+[7���\�ܶ��O���6��S�3��S5�:���/�ճ@��292�-�&��w{�R+��S�t�y	�� �E�ו0��q�<W�E�������~�+i�@�a=m����_��{�A`q��ǫ�������h�����N8=�wQ��tx}����J��\|0Xj�^�=�`4�Sl~��y��z^�ӯ�E�a�������T�=[���<��yZWx��*�\������~�w�N����xjB��'�Ѯ:?=A��^}x�#�l���_����O��S0p���.J��PF�]���{�ݝ�J�~[k+��/���ddP�C�'�L����!G߯d=y���$�lj�YB���I�T󼶴�	`6���'�q����8����D�m�?��~��b���;V�5��	��;ա(S�/����!\���}/�w?�h	6#��޴)��;��;>=�mN]�UG-���ʉ9�ڢ�3�Ӌ�"h���j+6 K�ۤ����"����	�Eu��A�q��N����IB�c��)��i�9�ɳ=K�����%�{#;E���;X�_^	���9W���`�gg��B�L ���/&>�q�&Ƽ�?Z�����gS7_��'�ď�)���T�/D;���w`�����xK��HU���T���<CNK(��L��&��X��]�AOӻk5M�V���WmT
t�ܪϨJ����й�����T:���HkGӬ(~�_k~��3b��h���m.+E���s%�dT��O�43Tb��P6��6u��@�hh�F3�}���|:s4u%�z<��%����߳<�!���gՏT��I.4�n�(Bl���k�����eBڟ^���5����Ok2>�>�=Lc9���:�{<r	�9��@Qe��/J�^Q��S+�~�l��jD���v% ��]?CvDj^)y�O-�	�o��m���by=+�Ga�}Y��gт;��V��B���Y�n��G�I���$�lԂ��kJ�l�Jձ�B�����g�_��i��iP��'&���w\�p$�#6o��.�	bcn<L���Q��#*x�y�8%�)ԇ���0gu�c=��N��BT�?��k��'�Y��)������m����U:�!q�3��83�C.;���ʁ�-քא�2���5���o�%�Jo��jM�jU֨�l w.���*��}��6�w�xu>է�i _��� ��3��K���y�����|�h>�߷��Z6S��/�o*M��1�e���{���k�MAy6_z�f�iޅ�U:���B��Vb���S�C�3/� f�nH�)��5k��)6���f� ���-�wYZB*�L�r�;�Z����Cq-_Nϧ����8��bkc-Z�����It�Sϟ"@����
~yig��e�C�$okU՚�>���<�GX�N兌�g������l�P*ۿg��M��8t�0z>*��LL��}��/��`�i��m���z�jb��\�b��T�
�;&�<�L�k>te��`O�j���W5������	1��}}����XK�U8wۮ^�R���O�71�h۟	)k���.'��>�7=�3�;x������1�HR�	��T�C��A����%��"O�8_Q���ܥ��}V�E�K$a�e�"}������C���#�͠�'��}bȂ���u���?r����J���t/U1:�;U
oOs���{���BFX�h(��bN�;*�\�ٗU��dG�,eW���p��~�����s|��_�8Mk���e����S��	��\?���^ȩ����f9��H���]� Cֹڿ�+�ήQ�Xb�K?.s�����0Ȑ��]���ޒ�}{.�dۏ|�Q�S�G~�tV�j�͌Cp2��c���y��(�Ř� �ڬ��� {ʠ$Ӎ~�Z���.,J�$4�f�-~�b��̡�>^�;ű`�k�oN�ث�Œ�⒏�������w*N�m���m�#��lʏ,#F�g�2�Ǐ)�~8f+�!m<A�� �"� ̂�����8������d�q� O����{k����Wq��H��GUG��=d3)�h񬚼���q,�������W�1��M:)�A_EZE}**(����"kqS~�gq�Jh�T�����[��g�{�wZe�����!�>�e9��[s�Q�ld��:�᧪=��S|n���˦uc��+��������@��@P̺B���'�[���.
��}�GO�F�Vl	N�&��uw�;&`����y���$^G����Y�1�|�l�ʤ��Q.��i�}�|���6x�I#KJ�����<�!���:�,&)�Hb�]+Y��������}�3NRj� <�H���"�]<\���Uc����j�Z����+ӳ�a��IߐaІ���PX&\DL/�#D
�=��Qj��"F)��d
�X΀�S&U�e���{�a�UH�	��g��]��ܟt3X�Ɉ�~�+�I.�v4���m�,�d? ��h��q�iܼp��}�E�a��P���<D&U:Q_�,Bd7I�HqR����b�)ǎĤ3V'�G&��c�':'}��2��^*�m�I�$�	%zB��n�YR��5���?��&��E-���*�cJp�+����1��	���/��r��ȺW�������"$aoʪ:p<�G��C�̹°�ʼ�P�G]�-'�t���T?%Q��j�ξ��7b�vzI�b%:�	�ǣ� �X7���?g>�
����Io�#i�-��hlZm:��״T(�\��>�&������:t���iw²�\;�Y�L虢��I��q?]5O| k��!�m\��f
����4��f�`-�!�ڥ�~\���Pٽ�R����KMc�S=r#�2���-Cxv�z5�'�Nr����;����ŝ��O�޹&�bt��������]�^������(�f�M��Ƕ>3^�{ejv��l���.��29�U3�������X��ȧ�棐�3b�e }��nv4j��e�A�o���_�{8�?m5m��;Ԁ�G}�g�؄����:�_�=<���ۍ��$�#D�E�~1�)�l���щz��h�08��.N��JZ��u_� �RU���K�oa�V݁�x6�\����*�����	ʻ�0�-Ԓ�`E�UMI&����NB�O9�<�?���\0|I#��$��Π<q�,�uOƖ��6��D�Jx��6�3�]96����:�..�6�Ȏ�n��`���&ݲYg	����7��e+3�g����g����l�ߞh!B$j3��څ;)����f�����@a�d˗jڗ�kmf(�:�iI��ЭO�[��M����2oOs�Kj�u,K3�O����E�cW��J����P�3�wT���]Ӓ����dn��<�e��ۨ߆{��H��B�W������G����\�>V�'W��B,�L�����q�MV���%]�[c����y�J6M�o,����bO�PTb�^�oSiT���#/Ū���J�,޽{D+�Aרƹ)��Qa/��\9�+�s"V�,D�x~�D��og�æ~�ϒᡎ���%�����.�Gnӑd�+C�^�`�~x�{O��RU�m��-U���Ƃ��+�Ű{��$�nb���п	b�,��}��f2 j<�e ߌ\���oQ�l;:�-.3�q���	͟	��W%w��ozߦ�C�̇�_��$H��|�q埠���؝1� g�����_C�C�W���P"1��]�Qy@N�k+�P��~�[T�ע��W�I���Z^�u����pz۷��]��X��fƷD�<�k�����+��'|ɽ�|[$���W�5�onY=ۻh�(���O����������"�E��$�'���X�vg���?h�e��!0GDW���rG����W���~�h��XR�T�/iĐ�"��{C�I��~�Le���ꖌ�w�$�޴��+����z����YI_�=7=���S+B�õ!�/�C������Ӷ@X$U΄���I����Y�=c����R��J�f��魆����uG��3J�y������zOlm�s�R�8�Y�yT,��Ke�x��e+U�͑j�M������Z]G�����el�����T����1A�g����"��剨���o.���U��
�qV>���(�d�通	Sn;�:_�dRG*f�/�q3��F�e|�(����i��C������8�d�!^1��~-����<A��E��ad��Y?q��QV5��g�ox�����s���`���	<�|�ŷ&�UX�����20�0B1��8�p�p�/F�c}Mnq�D^��u¸2��X�v��-�V���9Ղ�4��H�>�c�4)vY���`����@Ȉwq ��ɵT)3����ә�ߥ��P��^���Ũ�\�e[��ߋQy�<� ?��ߡ��U'�v6W8�J-f͖���D--$��d�z"����@�{=��k;ͻ�1������)Zұ$�+�-����q��\����ױ7�A�{�p|ģ�,}��jJ��}��Ā���a��v�?Χ�S����C�U6�%_��}𬈃�m���"��,�P�щ&����ر �����(3c3*�I��5���έ���C��Â}lpk2�$��9[��꓇ $R�� �+�P���畂S��Մ�YQ�uN�aKcħr�x80��⬷�5#�a��l�M䗋�?���^������d;�i/#�j哤M3�����OG�P�h��+Nבqb�x�����20�<�`m-�j����Ef"�����H�z�$���5-D>�?��Y�����~}�Rk롺H����MP�
��|��}�t	(�:���ʍ:e?̰q����9U�b�R�V}���;%u��?��7�h:��҂��+�k�F���gl��7��5�����U�������f���,.�}NܐS�-���g{�N���7���J���4~>���uʼ�
H
�Y;g՟�d�>p���j���vz�q�o��-�:Eu!���i��w���#3��9\�f�E��yEzYw��]<�o��|����_C�
���ݷ�
+�T��2OK!$���&�[~���hT�ߎ���<�_n+��J�ǁ��֩�4O�kF������.q�7��k��F�W�|�
��Ē�2�|De�|�Q+h��g�����u4U��{�9>��8�}BQ�_-�[퓐��S���"�k�O�=���~5]|�������ͭ@�E�-�c'���q�'��ء:���U�H�%�N�K4'p�쯐R��y�����Ok-HKŗi/�^K$ǩ��2�J|����-!z��\	~���h�������:1A1̶҅&�!W7��� ce鲓F��Z���"aI�ڭA���;e��8V|�r�-�3��ew�٨kp�k�Q1쌤�lNg�q�%H��:������/�{�M�+�#��x��Ά��l
�g"�o+��wnY��N�k������[ϳ��#`���c��w[��ٶ��`)�V����a�0��V�����#��Z�ܕ��i�S�ş�纎� �]� �<���������.�n̦�f��Ǒ�㥈=�)� ���#~hks�9#�bc�/�x4�w��2�*Y�w���G���Q�sȟ�ن-���6���9�\ne#P*!�EhL�Q�=ƥ\�I��� �+`������*`J��%��"U��S��w@�.D.�F�ܥ�y������c��;pid�
i�٬��Dv�5P����K�N"]�K��2�]r�bNS��L�+Dh��p�fw���Đ�����'y�[q����@9�����2���0�pco�v���L-�z�_ʭ��G�`A�§Z�J�`N^�����~��3�y7�K`1���$ŏ2p=I���h��X�tW�LACD�8�m���]
�3�.�d;������y��'h��bk�`P�ϴSVx�l���L�f��c�o���[�,��ґHdMa�j~�~��$Z���_��ۓCp����hi2��&�B����͖�D�wP��i��Æa3G�+s�v����7���E��:����k`��M����^ǻ�m7�뚅�o��)�7������
11'P��z +����?��9�L���s�M�H?֟�����&q�V��v3�;t�
�:X�����< u��2�2����4�Ң_2�	���i{"��˂v��&5k �W���&���ިJ����2L�A2�>���3��r���h0���5�D�Q#]��p���A���&���a�������=Ol��(�'6�@�&��ލ�=�9�^���9� l�ӸrC4�7pG���i����#��SZ�u��YwP�{��-�21�QDŝ�\���_	����	�o3���ÿ.�Y}ܓ�,����A���JA����SLNe؉�5r�X�o ��� �Oa��x�9��Ⴧ��K��|O��M`@�tQ����4�֪��h�
_Lӊ,�/�s�P���!,�⺛A]�M8���T��88�*��\G�!�	u"a�����~�c@��������0�@�l6�L>d���קT����#���ڸ�[��Y�K�K��u䶱��dӺ�Q
o3V@�r/������=^j�w�{ee�v�j�4�0ZC�k����>�'[T��d�Z��Va�D�W	��U���
��J�� ���W>�(��]������<�7�K@�6-��R�&C�G���*AC�=�(>'7�ɸ	�A�-L��U�f����CT�|��¸�cKn�${Y���T�f��5F [�����	����4��=�x�WV�|ٽ�{��UFܭ�������q�7�1�Ď��,3)����g�������n�g���ۤ� ��}����J���d��?��D�F�̷3~�4�䷄cfV؄zGDv���]�'������6�o��U��Z������u�o��Я�uͳ5��e��
r];���]�P���`�?�vwU��'\;u�����f� �^X��7���,��I���vOL4�n����Dǚu3��k���~�f׹�~u�P�g����|�J�2~�Hy���WfwCC���e��#��+�����ˮf>R�դ_�$�lOU��P}��W����I����$��u9��Ԟ�p+ǈ1����,)Tޢ�)�Em^�����!�fK�H�zVgY�V�o�:L���(� ��g,8���y�ʺjQ��׻v�4���Y�r	���m
�j���b���ӉB��9��CRV��g���h�@c������������!~���r՘8~#��m�e�����u~�S5!8ɣ�E�������j�g��|;�hWN}���	~UJ}����ځʣ?v�9�Wa��$�������S\�;���h��!ImE��;���cI��޵K ���S��l��+Y�2��6�Y�W��` 5q�������+ՅST2D��\�V�f=�N'���"��/R_x��ROwL	^xB�VĀ���@U�Y��|QM�֒X�𪍆�����o�H˸���������@!h�.�&�������	;'��0�C-�Z����r	���������%~	�\C�ذP!�'�x��ąSxcc�5��u?X`="�p���1�N�J�R��;�h��av	�����X}������@�2'�["�i�P��˟V��z:ɉ�N��E_�҉��"��q�%�z��h����i���!,{-���dK�c$N�J�;�|h"�}�Z�yT�9��7�U$,t�K��˝�����[�)�t��<.�.Y21n��*I�н�W�sZ�1�:�==ی�@�Y�P
(v澃��mr*��OK�,{��15�攏~�ׯ�j���c�gj���9hCDT�P'���A�QV�M���o�y�Ǽk��aV�8I� ��_؞�G��U_����E9���>�h��-�%Y��7�=� �g��e�9��V�B�/p��ƞ
�<{Dz�<%�T�@��Ӊ�^ݣ��v��ٔ����Z�?��a�&L����ۯ.573�5��=����N+)��Iâ��������f��������CB�T�]�v��X���&�>'��v�������z���,������w��'!�_$C'�b�&��A�Y����8�b��e�(s���u��֥������I�4��F/��	bD.;�KjL<��Njk��)�E�B���J��-�K����::E��g��	�25/�ٯ����SQ����/k�kli*�@Z�^�r��=u�|+��t���qU�3�x��K:T��j�� �5g)W�HH�b���w�<x���� ��;��Q�wǿ����P*��+I�����z�S������M�4��my���L��+�aIux]|S��os�fX�B����I�=�~�Mf������P�*�Q�$EX�F���?�*r����>T����Ď����D��u=a�0Ƅ_9��1�X��I0��Cy�<��.�Q��%0$:ZW��D�'�v X�����>`�C��G��|V$�0�~Tb���#M�.��-4� �2g+��=7�+����� �է_q57E[kt�9��7{�n�܁�rd`9J�)S�ό���_���C�$�9ԥ���4��3�����Epb�#Od�E.���ѧ[��Vz�ؘ0��Xw��?�#�mO+� �n��L�y��� §U�5�-���#6*��:�ȣ�t�^��,+�ۇ%�k�!���K�	"W(T�	lƯ!�:���$��!I>Ş�#*�[m,��E��rVy`H �	:K�ξM�+�v{���c�����w��`f{q���!�Z�$��*�W��"�?��l���Dv5yr	@H�NAK0�%(��\�<lV.�}By�q�wE��,��W�ض<jj1�|������'@��SF
7���C�}�F�M��\]�kkexf��҇f���#%�/Y���&�n�\w�������u1[�: ςqH,��D8-������oxGhE�髤�ۺ��$=���g.�|rޅ���u?@ܭ
�mz�C��Į��v������[�l"	�q=o���V�Y�kŝC�X�TgJ��+~&՟ ʡ�r�! �W�7�J�����s�;�ߌ93^�h2]����l0㞬���љ芞|c��6����5/�8C�M�a&��<U�K�l8N��fk����Ϥk�E�_U&ʢ�a���>˞\�̓�g�ŤY��aG�}r�:z�G�-tBr�A0�y�T�z W��Hl�x������2�_�hi�#�60K�yi�*����u�����ɶ�xʉ��d���=Y�[۟&h�IE����)����������"�&LT
}�+�Ε
ݳK��fy�{c�0�8y\��.��w~�Y=�0����c�щ?�7��d��<�p	�T�?��T-��pL�������OT8�pj�V-.�wT�Sq�
S|��C�1���S���;i�N!hr�z�r$bio��$��_��K�r	XMע�rPVl��ck�3�]_�QE(�{*���Et'A��n�<-���6��V��n�8�����y�&GŌ׻9�O��/���>%|�*I��h���.��-��
�r��\Z�иV���������2�*�DU��GOؔO�����8��������/�xN���z� ���QhѨ)!���b}-��ߠ�5�Z��yC�|�\�r~���ng����=����$k.;E�RC}�h`̤�j1/G�����]���g�z�3���4�/�g�C���5�>�7)�a���?A��g)�߼��֒�K��f��{"H��Ag���Y�o&H[���;s�3�̰!�ۭQ+&щ���W�/�z�����D�Aw^D��h����Ťc�~��@�d4b�����������>�A�B9[���f���]���.\���^�H�I�K-�%�a�{m��2H{���h���%`�~��?�g�k;X�>�&
�"�6��`��5��R�lK�^e6Ð�iA̼��؋,�ݫ���A��m����L�l�<tՆ���5qA��X7`�Hԟȑ�_*��e��9��t�
�ԉ��r��*䶵_�けl��n��؆�Ql��%��/r:3���0�r�@�Ld�M��	s+d�Pr��Y
�B��7]`�'��3����&9Wt�3$������1�B���;���>�ɋ�=��;���q�lٟ.9�
����(���<8X8xq��wJ��^S�I���ҒpU��NG$I9�<�Ѿ�~&�T�g��;��2��/����]�M����}Ņ�O��P�M*�. c�E��=��1M�>A���h����b-{K[�����ʮ&�\� c�/@�3��_�!\��D���_�5��M�n��	|w$/ǻ)	?@L�T'��}į9od�}��֐ �����R5ie�a�����"�i(���ʤ���s_��[�oX%��P�FB8�e�������L�G���o���kcMs�m��B(�E�]e*���~sϻ��S	\ʾ�`��P��~"��ƭ�:���,2�r�<��lW��ȸ6��׺j�Ǡq����R1G���xwh�M�yy�&a^^�7�
��s��;�)MC�m���S5��b�ȼyU٦v�m߽ﻛ�m�N�����eB�������s^r��7�d^ԏ�?Sc��A}f2ª������R?ؔ{L��m��@q�B�Gz �m�5ؾh���l�����q��*��~-������R�)�mc�s��LFnL~)��R.��	�7�Y����<�eRvu�u.��T�\��ȁ&���D}�{h_$j�%�KMgS��&�[;f��q]��s�X�B=�7�%��WFa��ϫ����L1��F�z�&C\��M1Ik�c[G_���:@�Б��.�TD��������nw��� ��N�G�f�䤒܇5`sd!�e2�a1�^%p����wq������ v���ZZ�xOi;�"W�:�;�}��Z�׃���J���Y?�IҲ����(ڗ1����}�9 �����~�����UK �^� ���8�0���D�N�Ɩ�o7f)O0w�����`���
�PW��d�z�C�� �k�Lh2N��'�Q3w�&.�6�_.��$��2�=�9���r��%v{����R�E��ҍW�>��#�^?5�T��C�Z�K�΄�x��������:��/��TR�.�n�Ή()��ftJwm*�% ��T�A:G��nݰ������}���9�������{���Ԟ=��-]�(H��e��y_��}S�J�?k�������qS�1�O�޲Cͬ]��;�EC���9X���l���դD6�$�]e�;��!|�A���"g��k�(k�
����T�r�f�z��랢7j��o��&��v{�ծ?��*i��Q~�)b�S�I���L�A�@����Z�VR�����<5�n<�3�q�
��"�=p��~��~77i٧��4��7�o��t�.�T�Ly�V4��`�|q0�����g%�r����Fizu�7�f$3�t|��K�_��D�sٗ��cQ2�[���`���a�����k�baJ�ҽ����R9��7��r��sy�W���t�=+۪8�ӌ�3�8��N��Q^�����Ђ^}�F��$J��i��;��퓤�����eM��Ύ��۱��HW�\����f޸��G�#��qlz�ac�������ν�7rs���w��򔻐��BwN>��WBt1e�h6`��6m#�^�Уt�����Rؗ�!L^�@����1�M�F��Ѫ�Q�T�ٍ��캳<ݏݻ�(�\�3�������dE��UA�y�.>��oS�ЩFuM�˰�8��\_��5r+0��Q��6����+0�)9�O���G^���_���֒9@mF"Țe�emH:�/�a3��s�he<��S5����������(۾�Sn���h���#���|�Z0Ԅ�b/ ��F���	1��S =��f�_-�ya4�9�%�������#zgVƉ�l����k/�^�'�m|�E����М�ci�A2�n�>W!1_���׸W-^��Q�@�u���"���o�E�-P�������j{m&n�OG�k��ɝ�:�{U�Q�s7�ӂ>`��O�8�D�EzT��o����a��F�Ò��I!9���`��	��Ú>��|r��6�kh�{Ħ`ǐ�P��qf�2�P��?Gkh��]��etӪqh=+�)V�R}�U1@��6Z����=ō
`�
�ư�A��l65rw��B_tn��H����|R���6:�S�G}������g!q3�a�Յjh���ǳ� �Dk�<��)@RV�)�(���6�k��=xX��r��y�@��w�C�r�H��i������G��.q�."ڞbV�lb�ʙ��Q��F��cj��/�	���1(���Pj�/�Ux�>'8�^���1����]h�4�xb�vl5:o�!m '��<V�����5�$D�H1�iWݢ��W$���x:�ԑ�?����\����#?�� 2m΅�%#ot6�:e\Z����������-�����S�=�4;`H�*)s��{�{z:P�1N3����4+�N�/"����p�������� �����oJ�`u$��q�~w�~�$�j�ԸЊ���^�\��k���!���Ҫ �Ȼ):��SVe���N�O{��N_.z���E*0c\���D���H9�|G��y��
��[V�dU���>���2��9G搡�y\��ӗ?���O��� ��m�"9Q9L��j&��ֈ�*z��JM�^������8JH����5���QK�ɦ#ENU���������-�YJ|�|��a_k��T��<56��X����G�|~�O�Ȭ����7x��m�Bk/-�_���{r������v7@������4<��f�u^�m�ٗf��;�ᦄ�xF�/Y=2V{�d��|@��T@��B�p{�L�s��۷D��P���pHY�ش$���d�dF$�r+���&-֩v)� �X�j�ڵv0p�Ñ@EU������Fe4��'y��BW��'>�pj��9���1Q�{�����B�{�_nb���t+���U�I�ږ�����L�m��w:]�0`��۳���#��nsO�B6f����&��U���"sqݏ��E����o%�3���I�>�c�{Q1��i�v���T�?A���v����R.���)��FЍ)�������Q�|�t5N[[n1P�<�vq�j	�zRY��эm$x� ��f�Xj�޽�e�(lMW�U������0�k�]�����	�`[�Z�5�60���_�|��KIK�k}�Xf�U�,�v����1Y��(00��"����=w�PP���c ��#���Y&s���ߑ��=�Y�f��v�h�a5X��nVz4xp�lrr����9�v��a6^ݤ�BJ�R�bm���˛�[��+�ˍq[��hFq�>��)��JR�&W��6�=p�mz%c&�	oo��zVv�p���pWS��z��(o��X�*6��� ����l��(�#V��t~-j3-ϟ�s�x�)��߭�)�BB����;p�X�7RL�!�b�b�N��髀��uߋ̒܍�7\�ۭ�F���G
-��%�M�BM�:��T�2dh��Q���s��s[2^��ބC�g���2�1
�{
��zNL����)[̙�Mlt�x���o�o!�I�eQD�?�,�Z�Ȍ�lL�}�@]$	@\��+Υ	B�-��[$h.������ ���s���ZP�7l��l��!����j�vW��X�0)���cs��Д�"� '��u&�n�ފ�x�A��W/�9Bd�yO���0)'_�Y=�JS/2��D=�p$A���߻H��^|p���`�5�6@\�$+����?M)i��O���+�� K���_O������`� ˷%*g��tpd0]aǪ�T���Y���>u�{��%�y0�������ｸik��� P�x����.�bX�rDԡЃ�Dv)"'b)�н��KsB�n�_�6&��>�#�����'���;����j\+19ta�%�!2�//�V�Q�RJ���u���u� ' �x�P=���=�֎����,�k��Y^����|��f�Iw|��6�<x�I�E�Yѓ���uŉ_#4��;cR�?F�{��d��˦��"�To!D���z5�����Iv;�ؽS�_��ْ\�Bj]� ջ�}�Ft�rg�g���|_X�ݮN坘��
k��N�w*�h���'�DB�pW��$̒3���h���F���q�Ex���\<��S��x7ĩ'���^h���J��$��ay�"LP>��a�R�C��P@ ��uR*�u��g��T7�75Y2��)vV��nA�2w�I8�L�];������{���l�Z�u%�6��K��ݪ�P{�rt�`H��`N��q7�������+�\�!X�t?�#{y?�r8��{�����^�G�n�l��WWp����P�3�{y'͞���H��?���ܽUƤcO�pz���zU��������	�9��:��?!ox�I�[��[��c�
(���}�MEE�}HA�>�ϫM&���	B��3��8wK'_�1~AX�z�c������$ �J��eR�[t��>r���,�/C�L������ǻ��R���"ጟ�Ac�d�ngE�4 ��p󁴼h���=!bIy���y=]���t23����̪�.�1�ߠp,�b��U���.�ѽ��lD �Nϝaղ���dN�H�]�Bܧ�0@w3��
�*���w���]z�?�_�(Pae��Ҹy7P�}��l0�{�(e����\�sQ-��s�c'tj����W�/"�4v���������䶳��e��Is���/Mn�2�O�X�o��t5�Ni�v��y	�d�2���MBg�uWl�EV2W,d�y�4�K����_һ��5N���dW)��q��H�E���ӥ������9��$��"����x �	Eh�z��}a��:�yV��p�!�f!�ڴ|2�o�/�v9st���a��Ў|P ���G)�<(>��?��?����
fU2ƽ��ڈ�\b�fj�3�#���Q8��zC"B&��C�I��Lbp�������R{Y1$�@�{�|&~�����z< �K����
�6w:�E�-��6sfe���P�q��O��5?���*˘ĩu�jl��&eE���.5,��x|e�WJ&*'؏����Վh��O�އ;�5��qh\d}{������oF]�5�@f&�0��xfU�/��:)���W�AT#��%����?_�{z����a�2G�Pu�c��Ws�Խzd.������[���3_�҈�	��V�
�4�~�X��2.����b�dB��4�јm��@�ކ0��(��*�)�&qY&��e/�zt�����L���:m�We7�>~�����>Q�ӕ(�̯pB~Sl1�u>�e�t���r�Oi(f������>M����Gf�kvTEZ�-���Hi!�t��U�	���M���TtA���&f�AsG��}:PFڣ���P;��p�%C����vjэ�W�n1������ƀ��zg�-��aG��O�^;� �����oߥu~��@Vz�Z�N:�ú|0,n��<����ngj!<�q�g(D��>f�f�;"�(XP�y�lj���Sh(����_��<7�������A�����^�o�~~�K�K7n 5�O�h��욌仕�{}i��6q�=7F�T���+n���h~��ͩ�0{��1S�܂J�������M�z���w�r�"����V�iV$����B��ٲ�߽{.-ͱ�]{&��b��t��΂e���Q��T�w�/�04�v�b���I�o�����M"&�*���H>����P��1Ԕg	�O��"wR}��d!>�DXZ����bU���\�*�3y��og���D0�dL'�b�|��a���; X�j��O�ic:��%�hA���
����F4b��
���Ѧ\j�g6 #�?���K1�qǢ�kA��&�w�<��'���^4M����M]�-~u����[��cX���v��a�_c�~yJeNq������/���a)KU�C5ud����JD7��?I'.�c馸�4��.�v�C��U����+}2����M�a��2�/ԟ�}Z���
��`�R~:�&��ϥ�2�i4�>kj��x����h�ӗ�����j6�3�%���e�)//ۭ�=�䫗�g�4N� %��T&��9����O$���ɉ���)n��2�����]��護�얃k;a���lf8�/e�xC��.��@��{&�n��#B��ZN�y�TW����A��Z�l�g6���Q�82�`eΤ�4b�vB��/w�%��ԡ9m�7��O��}��:#�-U�"���F���T����g����ϊQ{�iF�N�����(��0}S͗h���#�����U~���_�C�w�^qb��b��->%��pi�1���E1>�^�݅���o�kƁZ΄�g�+��/|��59s<3C��L�ͰcV�t�m�
�)�mUʧtD��p�?���_d�y%�����H?��*kR86ms�>-�d���,��N��Z~�엗w|sA�ʟ�+��K����/��Ix�s�=C�1E'̈61$'�l�_�l��HVMf><������6V�;�������̏\���\�����鼴������O٥��n�Ӄ��Y�mv;�i�]N����S>�5,,fd]� �I��f�&�p}�F�Z��/��}Mۡw�*Z�������֡+^sUx��`<�b4�����:N�k���ҹ:�ܔ������U�� �w���\��h���B=��(�v\��h먉1�A���Ş6�-���fykp�Փ�Y��T��L��1�|�L�� �S���5/����E���{>������V �i�VH��Q┏tߘI�mE�u��]	_m~Ӹ�[�!ÁHM9{��B��dO��"�>.V�)�H,���55t��?�7�Ů6�i�W�z�Jm:;sD�]������m�:k�󽋧� ,����?�mγ�s��QOܺ1�G E/~��x�{��͕j���¡��ڠ��b�˷��A���@O�#��U{�"�b�ԁ�X�s8������h9��c��5p�rG�&�h���R��z�L��J'	�훻���%:!:�Xd���A@)Y��eՈk���Hh{����Tީ��ʩ��2���cim��_��C���S�ik#����7R�ݗ�̓�������c����3�2U��l����DKx'D�;	N�I����m'Ӏ�I�	>�䆱�Ӯ������:�{,��v����iW1�/{l�M�%�$�-�D��;�a5�nq�P�[��6�4���U؟lab�	R�,��<�L��0m#ɀO}�u����iђa�[k!���Qx�Qi_z�<�2%������{�.���r���էd)*���J��=�)��<
&�\A܍�̒����󿙨�7o�; Qo����-�9����%�?�&7��u����MC���E���6j�J���Ӝ��1zׅ�;0>�C���Ȇ�Y�8��z�A���n6���Y�a�d�dD0����M��A�zPm�@�Fm�}x)�A:�����Yjά�����"s�3��q��4$����\��WO����'`qf_�r�V�$τjߦ����l�(���d:�sP.��1QI�vX��cf�?ӆތȹ#P� �Sy!���/%/�]{j���,s6�Ҋ�Gf����_�_��G�T�h)���\���a�n��C+��kn�ٮf��ƕD���N����3) �)Wpt��L'<L��bb&k�����'Ϫ�5���e�I�E�l2+F�(=����TJ��z����/NNU�X>0���!3F�(!��ςʢ
�W��ʿo�~�?��[�잏�Q�9
ޙ�t�a" �)������ �d·Bt�	�]��ҿ�}��o��hn�����=l������<�k� �����M�~ߐͭo���iِ<��<���+�f<ٕ��݃��������;�R��$5qj&��ܪ��g�^��@��2�����Zb�X�]��"r���*s��;�W�������!���M����j�X˻��f|�=y���1i�����k�¹�7�%~x|'ܚI񜉵6���R['���6��'�H{.	{��c�@��;��W�t�	i�4}�}�l}���ő4��B�C�P����%�`�����h5���q��b<���wXi�򥎕Hq	�ˍ!��GR��D?��;*�4�և�doW����Ó�1�`�|��Ἅ�z�}�»�2�RW�:�2�7����e	ճ��y��~-�&a �cFx+�����q^��(oq��[@*��C�+�ÿѯs@����nt�}�A �M		XB����H$�&PMy�Xc�si�e�m�����<�L%�������� _��T��3�˻��rP��@�e�l���pB���|���ls'��h���%Lw7��O'ə�r�h]��O�}�t.o��e�4y�G�:�=�ac��e��sf��A�~�e��b�g���Ȍ����"��d���,�PF�M��5?�� ��ȥb�'���Y��<�S�SL� �c9*/)�O��-�;4|��f���WG����"����|NI��g)�ƀ��قo�>g�48�ղ��I�	7�qK9��:���J�\C�:� B�i=����T��>O���]
N�[,���~ʴ'h��bw�����}ZwّSVK����AZ���������]Aw�_�O����/���aɿ���}���:-=�ؖۺ��e[��,��N��_��l��� ��a�nk"j�sc� D����U��L�z�@�Z���oT9���f -�#*oJr��ا �u����>k���x�yM��M��1�C�E��_.u�*��A���ԭ�w*���<��v���kۣx��`�
{�+-�rJ�x�lf�5�c=H�����_�tZ4�m�C�
�d&��7�D6�S�4��o9��%.��$pz�I����%u<��E��l���K�3D�F����3��h�ąs�?̈́j�}2��k�M����h���.�vx�*{��zx��/��mx�3w��'�^�^h���H���!��R�G���<�AQ5&�7`��v��G���S\����%e�CoQ"�-�,l垞�/�8����>4S��5�'-X���}��ȩ��Y�	S�$����[�kQag����F����_.�R�����q�~�,[l9F��y�vN@QXUNln�A}���
yw���C�� 8�hNG�;����/��&?ļU�x�`�'Q/<�Y���MbFaJ��wae#/�o-��\��鵏�<M�cw��<z��=�R�!������Z��Z�TL%��_R�?J�}�y��%L��:���Bg�AQ��<���T�����c��H��X;���c�u9<����`�%��������9�V���_��W=��"S���kK9��!�ܼn�癦�s����*!O��k��ݣj
=0""����Q\�o�^Zͽ2]�^�+{s���<^�窠��|z=W1/��v��
L�zJz���o�{���`m�O���D�LZs�^>m_����Ŧ�aWx�J�C�rDW�3��k�-s<Lr���/a<и�v��	#��坤�5��;h}:	��KQ'�+/<@x�#<��];�r�:����&�
�=z���"<�{��n�`y�p+���-�j�A������ �'\���9t��߱ ��߶�A[��|LՈ��8�Q���7�D�F����2��0�Bu�8x,��*���H��9�s�>����Ǔm�̟�/�BV�Y�$Tg�u��^I���3�Qm�%���&�3�X��p�(�w�4�oI8����9�����b]�" �t�5Ժp�>�)q��f�;��<�.��-��;㲂����	���\�}�g@�ka�)��І�ou��^��֒:���鸩M��H7�A,�>�i#�����v���4��P�έ�$��z}��iL�LW~-KB�*m��N~v���g� r���sq$]�{�����m�a�2N~���@����ѳ�w�d�ɇ*��*=�%\W9ӹ"�[���vs������U�#v��gg�E����� ���Z°1���1�
*�ky�͑?(��;�� �5�z��j���iY��G^G&\_
B|0�ce��_� m�w��$���k^�
��9���W@�3a�V���4�0��t�/�ִͫ��G/��e=�/"?���1֎�0��p<�-�o_�������)K�do����,	,M��d�7؛��2�D��&/���1����(�s������0NwF�^֠����Wb�v*y�M�e�BT��!{�$"B��"��Ě�;�2:�I$��H����*��i7��L�GYm{<�7Xw1���"�W�5	Z�,ٯ�.�4]���y�VR[I$e�/��Wa&���x le$�U�9�#��N��!��nj��/|��_��*���<�.4ٔ����(�V�-'�����f��G�2^b%B�WlxW���S��`F�+�I-�]<�e�P���5�>���U`�堋UO�=&�^$ Pq+��w��� < <��0ݰv�L1�n#�֮cDJ������} ���8���	ײyynݯh��W�>r3S��U�9�5�֞��+�֕��QS��(�y�o�ϊ�rY���:�B�TG?�L�`����+Z�����]��Ճ�7gE�x ��G�����B��A+����Q�-�q6`A�����;i���PS�v<��r-0"X �AtR2��.�G/�Sww�ӯ^ Z����rx�t�F!�]c�oF�w��G�"V���l�qu٭C�:���*S������m�B�W;A�����	���;��L<���Y���=,@�K�b�TJ���[���_�&�Z��(<��/+}Iq�wE�~j�4F&�ӡ*ơȯ`��EfX�c`#��q2r�^�� ���j�)x�}z�\?��l��a��(�"����(Q,�  ��Q��94<.�x)ҕ��^��U�W�p�T�	�F�f�+��ܺޕM�K�+�W���L71x�34T���@y���Z$�D�"I-͚2��0����k^M����:¤K��hޮ~̥ǝ-"f�p_6*G�L���=������X�Lp�hm����W��#jU��N<�1�ٖ��D�<Fð��C���u���C��& ��KͿ��X^0X���!���sd&ezz[�}����*��L�H����h��?t�n�W��5�zh�A�HB������:3s;�s�?�����}-O��fc�Zl���1_��%���s���Ŕ�=��fI�����v�E^�P0�#�e�Q0���Tdq᫻c1�U�V�C^&0�dE��V6�D+�\� �α<�rP�át���#�����"��+�9[N9!��\�I�(�Ꙋ�"�o�9\��1а�{�{��-1ZK���^����j��o�F��?N�v���y�ue�e� 
�[!5{ku�N5x)����~�s��P�lXdP��e\��z����_H�0�_'�X�Ď\��M�)Y�  �\�G�E�г�y`_��@8�kD�P���e�X�X��|��oX���a�C ;6Z.�4�o�A�>V׶͞*�ۥ4�4.���`0�61��i�<Ӑ�,C��L�G�g�� 6�E'}���;e2�o�6c��uv���Jm[^��!3e��u����j=/�x^<��Z�{v�U�A#��*�Z�Y�bc�������k�W��eV�b�ngh�d��hn-z����)9KsڠC��R=��/|Nᙺ�f�,��S�e����`�w�<s�6�!��Y���4���˞;3��x��ޔX\�)w^2c��wzd'���E���m��ʈ@��v����4t�E(k诲���5K���9�^�"�3q��G �j�r�̏vL�А�q$De+����wk<h��S��"��p޶I�[����2]���P琥�x�q �z�E�=Kr��g���~�jR���0I�#���ըie�2�?�J\��w �=�ޱ��� �\+\=�߂���s��0H54�n����ص9�d�`�N��M6�&�c�u^L"���,���m�{q.2Zm�=/X�&hX�I<;+O���e{�q$EXP7
E�����l���ױ?bt��_�L��ƴ�4cQ9~�`�����W�;��L�i���Y�ߩp��Yo���t0}�^�TV[�/C5]u1Kn�pL��.	<\v"u���6��/�<AIR"��@f�1.�H���.�Ok��?��  � ���e4�_����~N<kv\3��@�
.eO���4�W)��Vm7g�ξ���j�d\��Ff�G��=�~]��L_B"�U�^��E���x�(�����n�I�|�A���RDm�ET͝m^mbyٙ��JvӢO�H��U�vb���UQ�����Aτ[���G��o|�C������}��/��f�`,�,ΰ?����W����L	���wt�~�#�_cO�ŷ=��P���L���T7�0pju�'L�V|�;�洟L�B#d�5Brv�2�4?a���t!��A�ū��~�o~�������������i{�l�~hɩ���ܮII]*�@|uy$!�nW�8�IV`K�
UĖ������Y��Ae���p�<}���4�Dh��|űԉfQ�ҧb�\��2�Y�_���6�#j<�X�M(����6�! ���y��8؍ڑOt��:}n{�y�?�N�"��iq*z����za���p?P"��E?�ԯ�D,`�L�q���Pk� g�y��Y�3@J��/6�%b=�w_6��$���J���6�����?Η�6j��3�v��ZB�Mؼ��FO��4x^KT���G*��q|v`���XA����
'.��Ez6?|��Ut���5E����G���8G<���p;�gkg��3�cKL4��v�y��	��ę�x/n�8�H�;���6�62��D�0�I�7��ga��w�[��dA�����U���k��c$����J �p���tc�?��'��9���vr�S�'�+���.ӕ����TaK~�q�+���r�P�u��Z� ������{��Q��}܋��B+�3UbKu�v�3�i^�m)@yj,��]�"��A�]b��>WƤ,��)����R�xF-/v�1��ӥ%�}���G�o��*h�-���RN�%�HT2�%�K�'�ۅ>%X�9.9Y0q�">|�6�`�#�f�!�:�Iq�v���0~�:=��{*�i�)_��Kt�hO��hdK�h5Q:�-�&x��Һ"�O���+�8S�?H�-w�<o��K��p��WC��O�P�9��k��4��$��k�j*{T�B�߬���]��h�俙��Ց����'u\�М�i���Xz# pb*��1���]�K�^<`O��',O�;����I��5����f�^D`�^��z�΋�'��������d��l��Ui�_�z~�+��c�O��k�,���"ϔ!��-'�Ͷ-²k�[3�L � u�?��&TV�����iԊ����:*z9 >�UʙTM��hz���V ���V?�>�����N`����7���}���>҈�1a� 	s��*�(��=�0	��˯GNWc�jt��Q�!�1}x^�5��g�u<`V���9�:��GΞg?���$e��	�3����9��b��LpNP\h.����"�ݲ��x�!�[cG��AAJ�B�t�N*�/P�t pQp�N%OhQIĉ`�
j�A!��R�����B�Ij��"�w����~��Cߍ��]����h'mсuٿ9��Z�/����c	/�ݒ�$x�j���k�%g��o.D���&	���rv���]Pt�U�;~�5����̼e�?��u\�����{7��ؙy�0ϝIL�e���}�m<�< �a��r�Rz�����ԧ\��y�b���e�	0W��m����E�)h%�X�R�����lPU���YDMn
V�#���w���z�)�*اMe�Y�tٝ���`<���ЖSw�Ɨc-9����kb��E���4D��-d$v3�@�[��Q��+ũ��w�v�Q󫼸��y�Z.p�[�{r
G���S���]��`s�ym��{���֚���Bvf9�(J�&H#~s��,#@a��:b'����T4KmO�l������ns�Л.�H�Q}�{w�ka�&l�$�u�,D�`�@�姎Z���Q��V��1���%�?(��ZA��ꉕ��Ď��0�9襴|	*Gځv�!�g�ʧc�
�(V���>4=��O;B��uC�n3֝��l�����u*��ȼؤ☋hX�����] #�)x��ǒk��U��E�S���B���0#i���$�6�<��ٹ�ea~t���oݨJ�q:lV���:x*0��&�e�PH�8��|�֍"�||�Q�����E���~�q@�WKdj�gk�L�G��<�)\{�c33bs$ϔ6gΌ�
�|�KR��k# �:�x d��0��C�"6]�aq�fs�vSF8�񴰽�H��M䡜oQ��]&�/R_ӟ%���;.]��(�]8�8�!'<{�kY�¼�)�a*�����ֻ����4w	���2of�i���F���>�q���5�$%��m�Z�'I�h����h8<$Ͷ��>|<1�Ѡݠo�:'��YA�b�\���ŝ��9���#
����v5LF~��(N�0:��^�� �(�~*+<�,6��ՔX�Z��ɡ]�uM�/Vq��>F�An߯�]�L��ɱ�Dd;��0%�S�V� ���a`�ڱ0b���)Ͱ���^Z����7��-T���G��΂��'�c����})d��;�!��1���V�d�����*���CıK�n:8��r�a3�K��~m}�rS뺟����A���{�V�|�/%��u���]�����BG=�ׂ�(���	��]�}2�\���&v���pOI���-+�}�����%�7"���a%����9��ѭ D�ou�&�f��� \��'�G�dtA�,�j�� �Z�M�*0#�p��LC�)�5q��0%����1&a�����4j�^��Ep�6V)�~dn�f[�kZ��=���0���.��(M\�����9pfVS�[�?g4��1*����O+� Yتu��+��\WT��o;R+V���Y#�kЇ�ٴC���|jy4����ѵ3���X4��|	�P�<��?���Ӿh��q�?q��zm�@�hU}Q��t)�>�3�� ����/��l#&����`D�R�bi@�X�7�$���m(��Q�������E�|�\(��3���ߧ�إ��w[��L�9����a�'����qO�N��F�ґb���Ml��.�Ȕ�4�8n}�}�f�>�7f�y�D��}�-x�!�"Ak"��xز�ikR\GƦ~6�X7	�(�u��@�E,�O�p_"�����W�u�!�
ʼ$��9�1Ĭ�r���=�;QZ�_p�^��"?ȿsr��7��8��������o��<�|��eO?Xl]�L��	�[e�7���t5e"�"��(`��y��?��"���Pʅ���n�m�D�C�W�E�ÿ�8�s�˪�
�9m��eC8ٯj(Xe��c�;1(7�E��򑵏h��]�����W�ث5���G�a������BO<@��K��;1w�v����L�vt����gr`}�Z�;�M��G:�R��x9%�m g#��`���@|�غ�n@�z�>L��Ε�7��ױ��V�k�E�C]���d�Pih��;=�D�u2�؂9�� H>�uӾ�)���ڨ.��u��|^#x~`��3$%j��rT��q(���w���`CHuH�4�Le�M�����߉mw���kx����w�m�;W�|���׈�P� ��DA�+�^������i��c��,���)U�z>�3���y����t��xCQU�R��|�g*RW�x �Y]����"�F�L[�A�8tO���]�.A�^�*r֗�����N���~�ig�.��r��f�4쭇�]c��4�oH�ݱc�3ۛ����NȜ�������˨���W��/W��֦X�5�YrΉ�J=.��R���M
��7z���H-���	eo�<x��\K�(�̍\��r�f�Zb]H�j��gF� ۙ;^m�¿���7o�6�i>B3\oSd��IOM!4ڽ�VF���ҽ�Z���G&�8���8��(�L� ���_m��ik��N1�Jw�q7|@ X}g��FN������n"����Sۇ�`V�ǎ*��9u]�C�-��]�}(ߑ[Ĵ�꿁 y_< -n,������h����E�6��<��=�:4���)8���l��FO���}��c����t���B�P��W���aV�~��/��f�|^Rv'���۽�8U�H!�Y�Mj5n6�F ��Yq�.\]�W��K=��Ȼ��?
d۟�en��9K�Ǭ��}`.�<�0j��	��<�k����̈́�:ʊ��jg��ۉ�x1���|\�{"��-k0�{-�p>���c]K�����3N��ۻ�M� ��*����K���q^��x@��"��ڶ+5B��&�]�R��˸�8NŕU<`�Ǯ���M�)��]_��Ly�I�j7��~r���%<��$�ʷ���R�t�^�*ݠ6	S}��Ob�tM�x�('�_��h<��}���W�4^�����8IS}�Pg���u�ߍx�weu�t�$Ne@�����)̵���JD5��{_u�%��j�P�Py͙�]�����-oj	&Z,>jE��(� Ʋ!a�5��R�q�'n~�W�ߵ��I̓��"-�|
�R�9پץ�R�1�^�IA11E�ɛ7�p×�WZ�_c#/=�v���%x3ɖz$���]ŻX�[�q���=�1����������J���5~�A�^���m6�m������k#��OM���IULg�n�#+ �g�wm�!%�Pw�GK���݉DҌHf��X-X-��w��hF����9<#��Տd@�{P��h���H±�Wt_2Y�ڭKfJ����+8���� PK   9�-ZE�U� z� /   images/8a9df60b-44ed-4a65-94c8-aaba687a6de8.png�{w ���?)�a�"{Ʃ�CH��ʖ�%�8$['e���Ief���9���{�����wo���x��y����|<_��	��P�:�t����J��}r	�I�r�������Gw=HHL�Hib�IH���(��z�b���荔���V�܎0���k���5��M��w�H�C:�wde0D>���Ag&����ܗC�ߑ��G�)j+^lM�׎�׺��蹡t)).)N���bK������k���k!�n����Sڙ�_�|��f����}�g'�����Ӿ��0����7�0��Y�P�Ǉ���~l��5��G޺E���|��6�֚��=r����""с}I�����Қ�l�7���������ϸ�ͥ�y��̗�}j�;FN������=�׮$d&�M$�.�)��Q�S�(����q3�C e�)����}�g4��K�)��>����K�s�Ӎ/"�
q���kk���g�>��OǁL�X�O�,���ٓ����;�*Mz�Ro~χ�U�<�e�A��8����T��N�e�չ?� �@ƦwB��'�c�K�<��9�C���<�tvE�T���[�e�-@�Ib��ΡX�8L�H��$�}<�9}��O��N�p!sF}o�ɽ���X������ �`r�GP'��e�c�>"�"�_�P4q�˃(Ҹ��jK���U��5��1��wo��l�.'9|�7a���I&�Dޖ�$6��ɟ���$7a����*�z{9�}M��a�E�߭�� w�q3�����!h��$�����?�*p�A���^f���^�>~J�'�܈%�%���0)|)��ւ���x���B,��`c"�'y��[�Q�M�M_������ƴ'!렝��[��+���{(Ϡ�����*�J(Jg�Wu7��e)�`��+����i��O��`��}��|J(A��H�F3P�H"Ƽ ��V���������E��G@~��_}���]Q�JÛk�]ؓP�Y+�/{��c�����*$%�H@*����O'%q�#���ѠXݚ��\����C�W]^>�x7���p��&�X=}�����`>�}��w��O܁��u/��qs��l�V{�a�!��}]�i���}۞��}r@�P$��w�X)�t>��g�WV��Fu�G�2>�~��/4��_��DL������g� �*�V���RQ�
m\egZ �gJ��P�����S� t'#|��9\�y� �OK�K�B�c�a<�m�P�&�7Z�1z��⛁nv��Ys���a. qA�g�"��u 3��8��~��&���������< �2M�	�:�T�0��ҧܟDz������Ǥ3�Q��x�OH�y;Z9���)��h������>xB���մ�������pcǡ���h���,!_D�`w�k��.4��L���$]&�ʡ+��j�V���*��"z&���nn<���Qu���CTq%��Y���
A8�8+SD��$�3W�m� 3�@�t�+��0�}�FϏ-nMs;M�U/J���Q��`�]R�U,��P�1��AiLMŹ=�<�Q=c�]�ߜѷx?A��j#�46��A{�l������)ϫ�v�AԥM���V5�f���^�}�1��_�\M4o�R�8~�&����窈4��a���~�)��ؕT�Y�1�T��	KVg��n�!'���V��S�����p6��B��	?��W�wLi+6%�a
?����A�e~�Z� уh�>��
�s�,�XE5�4�I��nM��β�E������-.���'A�e�{�~{�N|C�����Mj]�#�#E�����
=nwd\�N	k�;�J
c��6�bOS��G��!����*�Ċ���2y�D8*.��m�$~T��<琅.��Ѭu/��*�$}�rA�w?b"B}�o����ٓ�%��LʎS�����,Ll�	*��t`�a �? x3�#��*_��=�{�y�a;���qY}��ۛ��=��@��R�;��L�� ��������r�C���d7��Z$}�!I�q����>.�T�5�?+p���G��>$AS��]i�����s<Jm�-O�m�P�t�&]3�����r<��O�TG���6��i˵Ӗ��[�W��W��"���; w��yF�狛��{��1�fJ�gfR�7��=5X�g
��fhz�w�w�ϒ�A�Ep���q�/�]�i��!�Mmd���
��U:�߫!ߜ�(�O�ĨN"�'3�L\P���M�r'\Z�-a���h����9��f|U�`�Q1�ɵ�&dw	�}�?��/11���F��^�D��`�z���9x��?�П_%e��������a����v+3?����o��{��� _����)��'o=��c�{JS�rp9(���=�]$G�?ؠ��!�p�,� ����0�?�q�QC�����2}�l&��Eoܑ���&�b�uO�����(e�as�E�j�T�8㣎Q�&?��8��^��]^�9zt%΍(��S�o��,.�~K>SM�5QjzF��,�Lh8�H�SQ���{-��ּ�c,ۣ{	n�Q�c�^H�ut���aty�;�l_
Ū����퐵�j��0�� w-	'�}�/�� kv���l���Fm%N�e�e ���k@��(�|]:�=E:�;��Q��_1�Cp������� ؏^N���sF��sA�߼#h.��c N�����Z�s����v���S^q�:J�%�7��GSsd����S^��
x�7��߸��qE��JY4�PG4��/Ɯ_���L=��哆����p[:����0K�9xR�2�?�A8�������b�@H��;��K+c�!�0kC�!�ؔ:o5��\{���"�D�w�5m�-��׼;,_/l��<`k8�<_�������+>�+� 3�m2����]V��J��$�ZTq����j��X�nnh�}:�'�ED��'B�L�@���!ErA�P��~���*f|��Ĵ�)�0"��`�UA���'�9��DA�R����=�KSoT#K�Ur�M�I�`}tu���-�KL17'��&�al�>����R ?�����d���?cfquNٍ�Aك�$�ڋ�z��0f@�X��<RW�G�*�F�c0�+��a�%Ŀ�p=�K4�&	"&�(�A����BRؑ8GZ2��_�wf���oq�/&���)�D��g� ��R�}_^�����V%���-�,6��$��p6�H��6-���u4���{ru��ǖ��7��w�	��\�
O=�z��pI�Q���:�Hʫ|Q���Ʀ<,4ZJl�9�����:S�k�j�K�9������#v�}���BK4.D��8N8���!�u�Tw�H��
���L/��=f�����!��1Q��AB
-P�$v�>��՗��[�m��A7Y���MK��N��]8�:/ly��e$:�C�ܱ[KIUn��?d-ʭ�}�,�/#�!>�c�uWXI�:ӽ��WV�F7N�Y�A���x�Gj�,f��M.�M=�e�ː��lFv�E�8� hq�9?U�=E����<aYǌ��00ܪ��n���$C&p6AϮs��a����I���Nq8�*R���e���	�,��T�"�+7� �)��c�����Y�B�\��H1���^��k�[]y�6]a9��?�X�b�fM���n�(��J�N,�����F�m/<�v���:xq'8�◘�q�~A��F/J٤����y�5����[\2[�%_G#p9�f�>���Hd��8؄=HrW�_��1��?�]��Yő�6�H�G���^*�A���=����6�y7����U�o8ywd���z�'ո!�+ke��E`ѠVX��3��5�����Ӎ\�q�˟O�����u�IWs�Phjt��`��C��IO��;Y6|dr{�*ϝ-�ʰa���j��5ڍ�[�5�lTZ\��*[����N~~-*��7v!�'ƹ���	����[�"�,юU8+O����bs��j+�Ϳ�k� o�s��B�Zo�)-��˹{��
e�ќȏ�y�9-���O�jz���~u\�)�/�/��:�m���T�ޣ8�O�N?\��nذm��2�M�]��;LA�۶p�ve��P��$�#
u��Uҹ��x������@%�x#B�T:�Dv���r�����F°(��⁫-B,���2��5��u�ۛ�M?�$B�P��e����+�~��6:��
�5�!�ʥs���o����l���;B:w"Tӳ�])��5��:�MZ�8
��5���j�p�ѓ��!��3L�	U��ݠ�dSb0ҶMJ�'��%B�|�zr| �x�����:��*���4�;�
���t��x��bh�9�r��TT~l.��F�{��y�A{K��pm�3�7X،w�>+z6N�W��F��Y�Vג��-��*o~TK��a���^kwB� 0��@x�x�z�Q��sLժ�{p�;���E�_���6%^�!Ș�E'��0}�H�S�0����g����(�	��oJl�8�lv}�D�����-���?�KW�) �����~�P�_E/��$X�6)��0��9iisC!K��̂�t�ŬB�	�|�q1Gf�5�ܜ���ڸ߾�Fjl�ad�,��< �.��o[��~I�p}��apV;�7��p��9۬'Ɉ�O��xT�v�t7�שc�c�&��~k�-�^X]��k�:u:��}�>�e�rԲ><�E�+��	7&Y����^���G�C~�ЎT����re�2� ��׏�PnL}�x�D&���͵�T1�,�����P�zC��6�W|>q���)S���3�4e]%6_��SN�en\�l�)�Kd��l*���z�D��5��������_�pV��Ij�W��d^�na8{��"Θ[E" M��Ev��\����R�_�������Aم�vѭ�=<]U�s\��?���\A��ߚ_K3���O{y����v�L����Qп��x��E�R���u>�6U����5ί'N�.��}�#��%A��J[=Ϻ5�.���z���\A�K�_�3���@�,M��Ɖ���O Z��|X�{�M |����KFcL�P�eF2��b*���c�_(3�B����4kNe�_����ͽo���Ku:O̕���5�G�E[GS����P��!J-��5�V�k�������i�J���l�����$�a��B�n� Q���[m��a���t	�F��	�~{Q��^��|I�0��(@|o�WՊ0���0MfI�J��v^����q62�Ԝ	@�$2��|��~�:C��_	7Ev:��\ö�H+[����D���cYu�{><��pS�݉Ӽ��1ϝt��,��9��&ˏGu�	V�y�,��48�W�8�K\��WL����,��4�9�3��D��r��U�G!�-J;:�ӼIɔ����v�T}YU7�.��~������ ?�+c5�M7i��G����Q���˚�w��v�R1@����`p�O��0��v�5��)<���_��t��sf���;V������@�DH%�j�jLh�j?�4�&	q��E\d'�.�}
�/[���VL���k`��։�P��y��&Ll5�����Ɠ%��
�-wY�?:FN������Z*��뻁��<��g��:g��1X ��4w�>��.��۟�<n��v��#"�6`����1�B^t���s%Åz������f�|����X�¶`��<c�X����c�-Ya8�gY�b��M	��w�3z�f�sN������~f���	���x�'�e�2�l���ދ+��
���(R&B�~,�pfi��E
��	!�$���^2B��5:��r�U�͉���a��ng�=Vݫ���c#�ݸ|��L��D>�?�uH��Y���:[z��Z��wy ͊��ڋ��;�*���M
'��a< hʽ�u���H�Sx�]��w��&�h�F��@
h�w�~���fJ)��Om�>Y��.Ĝ@�S�nx����(����J����c�ڭSS�d�.LJ�dd��u�gP4*!��*�:ي�� E�Ge}"h��� >�--P����}�E�G�i�ȶ�����z��*]*�;D���NѸ7���p/�Q���8��WR)I��>k�}���>�	D���R�f��Јo��%�����)�@). �*kP��Ԋ��3�V�I�W}��>\����v�I��N#]-�s�4b,��8K$B7���{de��
[E�j�["��</s)�w����=w��=V-�ue�HO��MW93������aH�]�u�B"D�:�uibj�Y����jNfw�G�=����X�K����d�|�� X�s=�X�K�}�`�v8�μ[8�v��c�#�(��N��1��Ŀ�R{dCE`�<�0v)�C�{W8���qoѾp�%A�PW�*W�x7i��䉒NI��k�Br�[��� )v����y�<k���Mk���-IF��[/�G��]q���M�P��o����w��i������
�W�6���or���� �i�j���`�����ٷ�bÊ�'X�ѧ�+H����M�y#
�zfXA��'���D��� �vbǲ��1w"X�k���-�\w���w��B�Mk."���Ң�}�D�]DSV��؄��$'�P1�Vy��i�,׸�~�FWe�h��$�߂M]o�uk�ٹ�S#��|P �8�4��o~ u���vt��ޓ�0���$�פ@*l��`�AšB=5&l(zRGW�訄`dd`�Dey�:�{J�q�����eL.t����A}��_��t07Gmh�FAGg,�F�������"� 8Ϟ����Q�38�w��0�}@�^��P�����r5�G�|wǷ����:�����7z�R�<lY7�3�hت�����!6�T��ݗ�bǿ�R���53����-��E�b�޷�2nUKݯ`��!�%��<��?��d��A�2�w �e�x<g�""'!����A�<^�x�Ŷ��2-}��z=S�W��C��D��qm��h}A6c�6���^��H�ڛi�MʈN�D�St��{�3�\(�0^Z����Ů��X�U��"��ܼ��P����-�}d;�fʎ�^�ي����h^��u��)!�C��Nqz4Db������)�
h�-��U�/��q,����N�^v�<�?����P��\���K�F��K{0��bW����]7���a�o�C7�ߖ��e͋z@��œ����;���s>��-�sW;$l<�@l��u�l�MS �p������A<��,YG�jb?��:ĎA��U��������<�#�bi�|Gۢ1F& ]!����C���5��ڙ����7�z�� t�=f�h1�m�z��ބ�3���n�ڛ���F��^�ղ[�"Rۨ&?��i�]K&�z̮��i۫n3�ǌ�e���ul�F1�VBVW��lS }�Z��W��{ ��9��ƅ�t��(Mt��*]ewr������]S|ĝ�.�= ƨ���Bl̐d&	G���殜��F׮Q�4r���N�bE�"`~s�G�_%�3C�=i?����g$��k����o����]�(G\\8V9�\��_��ŉ�7�Z�"�m��&�W-�ι|�0�5q� 3,�i@<�I���x�öW����AH�͓'`�|
4�^��Q��ts��"�q�w����:˵\�b�d�x�`6=�Q���ǌ�a�%�sא$b��Q ?�m��1���Uf-���S�x`��q�cdA9�id�L�b�v�h��l,GUZ��ܼ,�(�����l���iI�Ԍ��p���E4�����d��t���6'�4n�� #�G�e)T}�������D�ݛ���Z��q�Ql�yݲ��V�)kp���Sx�=G�{�୸�3�N�������3�h�s��~PJ̧:As���;�UN�S�������?�,g�]�G���82]�Ǐx�\1c �z�˘�7���ސ���#�����b<�,���Ȗ����J���X�x~��&��&��6��-�`հ�P����Q���Z��Mkl�"E|y��c�t+q���؇E�I�t�|����-.��	#JA��nɔ;|�{��ڷ@E'JQ�U#L,�S���Z�_�d"����Jqd�2�Ӛ�DS���%ٯ�\��Ѿ�p�@���I*uu�=�[>�"��蔇���a��3����ߩ_��웞Y��a6-����1t�t�Run��}w�/֚��:L��."���z'U�g��0��"ݖ��k���#��1o�Þ�~���O3���:FH!�m��X�K�uތ٦f\\���]�VO[�EÏ��#Jb��~lO�]��>-C��}��ې�>����S� �Ϋ���q�ěC��/���Z��:���:�I�=w�x<����-�j�>��={"���0�x�����C����e�=c P^��@v�����8ȝD��$��ߑ���Y����M�5����t�+�Ӿ}���k�7m<sX]�2� ������wA�:Ouʖ��R�Q)qG�ƛ��Y;J�������a��\����GНw�%`��ƛ�� ln�/�LLR<��l������)���ӑ�%�RM]���.C���Se$\[�q*��Л�%4�?����y�$@�x���	�āV�8m���D\�����|���ؒ���?���7. [<5�D������.ʐ�U��Z�$+S�]��rŞ�!�}��z�/��&+ia�U��]5�8�j!Fg�:F�f ��5�M#�xW�3�]h��*!�OO�I\)��ת�)�i��þ_xn�BJ�������-P�˵�cQ����Ҟ��[.��
I��vw�Cɨ��S&���$��j�Pt�+����@+[;�T'�����Z����%;���#��O~Β�]/�����;�����ß�+5��O��7������92��+ȹS��B�4	9M"�x\�l{0#0K�!��2�U#����A�)��;��Њ
�W�������ʛ�6�k�`g'���-�φ�?e���u2���=�����4Y %��Nn�Eh�.��wHQ�&��\7��nu3z�xFSٸ)鲊�X἗s��?�Q�~E��
�9��IK?fː&E������#�������@�Q�^�H��+� �",����t��4+�\� ��Kp�]�;ؑ��>tkg������o�43j�u�1(ޓ�S��G������$�֡�|�4��$i �Mw��t�TRkf���]��-}�?U����
�g�o�w��~��������	s���G<�6ޭ�q~���+�E	�g���u���[��cxg��U= ��W�}is�))=kI���8��#�᳨9m<x�'Sr�6��D�M�#!��%��q��w�k�Gv|�~|���4-���"0&/g᭭Pf���׎�}y�Bs���T�*tup��T�,�=��~./ ���QJ���2-V��)S^�˕�'��_���x�ߣ��dw�?�R����R���3^T�ԩS�H�����}�?�gAe�@��C�/���/h<�s�+`Z�
�[~��3j�TY�=�e��F�� � ������MJ�;���Z�*��a��Ћ��mL:�z.�j��ݛDg���	���q��Y��0f�[�l[��<�"W�1����⿓��.|�����xL�[n�h��qc�_��	M9�e�z�W��F�V����]��tC�)�؏'g�,�w���)��*d�����n�s@��d�"/�p��w!k�	�,�l)j9{r���Ծ��*U�46��$��	�n�}2�B����� ������ĤӈXJ0	��-{N�w5��d�>�HE,����fLl�X�@���زa�ɗ�q�R��:�����A����#J����uj`/l��A~G�y�C���0��a�n�.���|��P�v��R%ؠ�L��7�u.W����Hb_ƚ��&�8ɆW��=|��RB(/1�0U�ޘJXLʎ;.�m�?����g"�J�ؠR����bs����ݾ�v�S�]+I5M��ő��� mG���v]�[�I��!����1x����6��VT�������$޷�����p�Nn�O#doE>5���S2���z�]h�����H���KtÐ��ty^�֌��K����}�� $��I���z���6��a�Ђ�Z�a��Ρp�9H�d�u ]�����>�OO!b�M��6'v],ǂ�o;8�u��O�*:,t��0���,�b5B@8�5�\{�:;Rl��m������y�o+�{���gg_�y!�m��Y�U��Ҟ�_���|x��1½�s���]V��2D���ևE��r#	�����-����m/��������+n�kꅎ7�'�ؙC?�p�&���nJ�Μ�7+��`q�^�9��/_s�Zc��^��iјz���H��	�w����Ȫ�΀X�@WZP5���j��e{�C��*9-N�te}���l��$��6}3�j�ߴj%p��|8b�7p�c����~]8!�m��Q��.��J�[7�7�*!��j���;dw8������W)˞��C��K�M/��z@�����)��^/�=�e��ռ,&E����a~T9��\�I��R�L�ь>�<j�N2/���N���/@�k��:�9����v�z�*�6�`iز�����\�p:��SQ���?v��������JvE�%�N�ۮ�6�G�j</E��Q���l**��j^:�0͍J��:d���Lu���ES	e��(�3˹]��8����r�Dɩ#��ݛ��^5R��>:"�ˋ���u� }��G���;���}d�J+�ӎ^\L]n���w��ݻS}����io ]"@%&ړ��ഷ��'�uZ�d��|��;z"__9XX�[�M��0>��0‏��kɻm�mb�z�N?��L5�er������ڭ��d{��+~bw:���`�A�5IL�j�a��M;�����i)�i�HU�~���VW^X\Z`w}�UVY�H�����3���S
�����w4�Q����#xcs�&u-_s��_�ۻ�8�~��2��[a�Ud^��`~ܐVe�p��G-�j��6�f�a#v�k�7e:Fxi4\Ӏmk+Z��6W��|���"���w.�A�'��4ŒȘ�]����AZȂ���K�,Gu
.>n�����GB�5i�T��	�����Zs��vs���AK��B�>!
��>r=��a/�b?c2��}n�eU������T����yc�z	{��ҭw��MK���s��B��c���R����H]Zս�;��¾�{h�<�O7�� +.x������m����Rr2ǝ̣G|��qv:қ�#�-��L����T�͊a�����辩��ˬjy�'��MW�O`�d�_u���Tސ9�:���Wtآ�p﹧��0D�im���S����	��K:L�)C��m��z������-ҩ�R�R�][u����J�K�H�~���J��ÌF��]�|]=_}gɐ,��2���K��ĉZ8X�"�HK�p{J0�Xw�9�ǣ����0�V��G;���t�����U�o��!9�����O�^�`�nsk<֨\���z��qĻ㾙�}`���q��Q�ѯ�q��Fo�W��Mq��ꥌ�ź�l��~������ns��*�� ��wJ͈cV�*S���"=�����D�ٜ�(|��%r����<D��%�G�&����8������K/x���_P�~x/=���@��G�a�����G��jʫ����~þz笚Kܬ��o�Kޔ�u�y�6�ͣ��6L�6M�q(U���\�&��k�A�n| ?@HM��2�= N]��#��7�Ĝ�E�)8�}k���O�q8����v��H��^<;���4:=�<�lf����Eo-��ý�X[h�'��G�W�Ȃu/f��
WL��>�VB�ӕ�^���/q��Q5�����2�W}�Vw0�Liqmz�h�j(:�x��%�M:5�[X_�
��ъ�Tz�FvX�k��>]����#Kj��)h�����$o>�����'���뎚%��l���&Ǜ}]'�r<�/�\���A���gk_�pRɡ"�ƻ~�I�6�4���x Q�4��J�hؔ� ��1�_�u?�a
��a�R�d�weۻ_߈�]��e�;�m`��V����^t�x�|6z�����:U��лh�չo0]�n�.4�w��ڜ���[�A��U����<���PU�6���vnN���)y��j"K�-ix���.*0U�t�M����Խp�f�NA��`�ϔcS�L�k���v��O��=U���K����$��-͜k�3�(��Y���[�/P�<$镠m�d����yRP��_qNQ���k6��x@6{A�"�Q���8GJۇ����L�b������Y����v_�_@<а����vu�z��Q���E}l�n��l����B��81u��V�m���9�Tzi_ǢJ�pT�}zf�`���螐�KF��JW�'�p�'Y��ۣ<��N�v�:��"�c���������Rj<M ��e��Wn)�f_$!2d�3V'�<���㚶�����h*3��ߖ�nO�ᶠ�s𫉐51��T�l
��q���b�m�ن7�ä�gM��U��X�ZUԂQ/�hz�\w�|Ui�7t����r�F�q��6��w���O~������>_�6[־���t��^������(��
R�o-|�[��@J�A6��HV���t��ٻͻq�e���q��(�Q��$�Ю^$uo*�V�6ŏ�]��'2I5�*fJ��W�g>T��z�GY}=OC������/q��ۗf\�ϤI1���߷�.�C�4O��}a�~H� h
��a�&����	���C������Yʸǖ�?�0V���`Ii�R@��-��o���Uf�TўYǝ�*��E����)���zDr�]~!\<�v��s���O<Yp����afW�*3d�fM��5VI�Nf�H:�e��U�J���舉� #��f�NvX��U>�U3zU�BF�iՇZǗ��(��e�Z�>}|��-�o䪽���*��z*�� l��g�8����;�Q�)�U�lTM'iߧ;ҷ��U��5��w]*CD�u)|
B�j-k��1,�n��T��Xp=y|M}����3;��|��P+X\I�[5�B�hRm@���͙�ugr�-a)���Rh3�9t��Y	�`�M	�6�ȵt�'|��J/�K��Z�!t��;�Ǽ@�ȕEM=vϻ���v�X'��ǲ�{�4�@9��KD<EEF�G��N䷗6��o�1���K��5܋�`���JG<6;�q(�:1C���/��5�a�Ó+�i��wYA�%c�no��f���X���+l_X��KK/I&��u�U��q����p�|4��4�.�昉F�`�=��
���2����\86��|�G6�Jj��vl��4i�p�n��W ���s&B�س�����G}l��n�O�3f^+��A�R`g�`���u(y�!*]Vж���):�AR5����E(�Jò4��#�n���Ne�����DL��d7�w\�<���ᠦ�מ=�n�J}�A��w�ѠB�8�ɣGf���q �/E�v�n�A{ͫu�PʠX�����c�B��@�� V��AVun�Ѩ�����J+ߎt��!,�p����(������<�Y���x�L&�Ny�]irٛ0��U�e��6�I�~�-�ϢU[��}�7���N�����	y��p�*�a抉:�;�4J]�@�m�E1�#��o���-���~o4��,�$^�.�� yǁX|���Z��J��3��]{���&��U�n����L��A�C��/�r����+�d"e @���>e�8���E3�� �F�[��y_ׁ!�R�n�w3�����ݾ�va�k���M�;�h��s�%�]x�OE�#2�?]q�I�OT:P��fc�zk=¹
ϼ;�|�����]�7\>�
�X��/�h�C"��A���8W�hVP��'�U������ߗ�9��7..��#�g��,=��v��B�_옑x��9Q��;|`Ag<Ȳ{��]�����������Uμ/Y�;d����Y�/Ç��[��t'?)�F�.����,�=A���vQ�(w���mY<��-��U�T����g9�K��gEe�.�n}'���}��@Uٳ��Joߐ�Ϯ`34���k����Z(���h9ߏ�7j5X��.����d�}h$�i5��U.���W�TWrC���Yc�	K�X��̈́ơۑi��^9��j�����єݕ���`t\Ѽ�����G���ap����^BJ�&�.�u�y��0�3���]dz%J^�����r�R�"J���ZmN�]5:�ʃ�,����[�{����l \tDm��U�m*J�l��XȎ�&0����w�����|f!��T�v�ڶ���J�Uƽ�g���� E����nx�M�pm����SvVQu~Pf2��8��4����=G���}��j�����z_e��L��%Л%0��Q�Fu�o?�S�N�^Xe��+u�B�P��������Nz=�N��)8�q�wO�H?��u'����Ņ�=������'�l�ᦃ���֬�

�ɇ��B����ڣ"��#^֟ڱ[Q�|��u�����roH�F��?�L�>� Q����!��1<��}����`Z��N�x�G�����U�mM!�;v�ݜ'ZdC� �i~-����M��.=S���e �n>���ǿ{��Bud`��B�B\��:�l���cu�ϔ.78�P�˅d��5��ie�[aZē	����}TlF�;٨�5F�'.,��ڃ��8~;�GUkdkSg\KF�u��	�����t�(0VmŎ�Ixz���g)�Y�{k��N��S$/�J-�����M��������v_�^r����a���b~nB Q�k���	8Ry���m�_��V(85AmPr��5#�]��'�;��*x��%A��`w��7�C7+�~$d�ËF�72<����50�1c�Ϻwp=Q�9��ϧOb��F�G5Q�=y� �_q�26�m9�4��������.� �qYj�E�G~�/t��\oi�_ԄU���mo?���x�!a��A`��ň>�P�b�~A�*#װ�Cn��J��z��ʏjqs�R�!��� ���H�xb����>�3#:���<�4aB;�t�_�H '�8X�60v������hl�Fć4_C�te�ޯ3(��	m�M��L:�q�ۙ�(y^�t�� z��2@��@�I'��6Sz����yP���U�-��^���Q�򣞫�Ё�?�l1��3�:����<���V��D���b�ؿML�zI���;d�g�wlr}��|_�׉�{¹���W̠���'�ss��F*��̈́��U���[���Ef�RW�_D��쫟F��S��~)���=�$V����붧��M�zf����PŅe1�"�Z9k����&hadu�Dt��]Q�Y�=�[<��m��I��z�۞<��)��e��o�R���iMTN�@��@�jPj�S��r�Y��F�����ee���o�7�-a��,�T�߉~�d¡he���"���Z�bp����%�	G=>�h.�L^yE�-q Q�"]~����]���v%P%�չ�r��0�Ljqu�)��+�W�9d���ED��QuqKt
X��c�K�#A����|�0V�z����k���B��W��&-�{_9«������ě���Y��c���8��O�
��g���\�$��.>�y��j�z��I[H/J =���a��)*���k�1cU��V뵖ڃ���Oқ���K1@�7���Vøx�k����߇.�cد`;ۧn%r���������䍽�a�G����'��a����&̂Qa�8{�VH�h~lL�~�Ž�S�2p4e|��1�&T8/�5-[wS�p�G�i)��֘H*ȱvm�Zp�E��͹�qz�����e�+t�YJ�����խs���#
tZ'�+ZCN	G��6p�{�f��wZ$�M�����A�V����_g@�ڢHԿ���z4��,�u�_��Ŭ-)�u����!�0�{�4{K���Q��Q�Y���h-�V弦�+a�LLD�����R`qIz?��/�Gi��НCL������فk䁌����V>,�;��*(��"�~����|��~LuY՞r�8�ve�\�tQȐe����6�P_�S�1�kܓv�T���͝5Q�s�d!E`W-�A�YQ�=���L]�Տ�w}�����&�Ѣ��4+��!���S/�h��s֏^���a�H�/�Ou:QsK$�3����E�7Y�N���8����ו�45��	�R�-Ԍ����,�!�M� �e_� 3����o��pY�оY�O��@���)2����P�-���S|a�H�b\�8F������e��3�SS�ò��K�ϧEit�8~�ys�q(��8��r_|.Ǘ�*F�۝������l�f�ӕ�fL;3��������	n��E����RZ����d%��4����3C��'o��n����K���uM��f��s	���zӾ�Q�Ekn�1�ؼ��.���za��~p\�C���:�}�4�;��!QH-�t�Ad��,�F�_8Z4�螻���1t��]So��e��r��;�1�p,chȾb�X)˔���S�������#�f!����v�q����ӷ;���Y� N���gԼ����.͸��x֫I�]v����^B�����t��lg��~O1�8R��Ȼ̆D���.w�wp/�\ӠIZ|�v�����y2����(q��r�����R2r��Og���[��?&n�������� %s�:u�9k�Zi�+��-�:ҟ�0��4��F<d�
7C|��ߪ�����/�'/�����ߌ�B�*0����;\��6g��Q�X�]��0�0������Y�����O�@�c|�G�v@�t{��㲦�G�+����.����4�$%<�{J֧T���J������q�dک���2&P���$�L���.Wz��݉4�͢��}w<���!렒}i��G"E���W�8q��-dg����,㐽��9�98��>�;��y=���G��u]��{|����Cy�G�AYC��� $�x,q#�8v����E!�t�.AK�N*�/)pz��X�[��{6_�p�M�
$��p�n���ҹ�J�?�>P>U'�-�0�z�;M{�W+(Qc*d�-�@������r~E��*�b��a�� g�O"N~Nn�U����<K�*ፄ##
O�Λ��_�Y%N��]���v�Y�EIM�s�ƺ�����B�xb!��k�K��"�g��c��c,
��<�M��&��{�jK�*���ֹ�=��t���֐^�c:��NZr�����!O���K��OY���������˳�>��U�j����'��s[2�ǾV�gm�MӢ��4N�%�\��tCt�X�PQS���i����h6B�b�c�]�1WY���1�j��Јb�7<ϕ.�	�Ppi�C��of�XW��%�h�h��η���7�qX�����Q*��<�/���v9D�-��	n���r	��=�A��>@�7���ڮ��gR��`�1�S�o�T���*x�$��a�����vHQVK>-qHF�u�4�W�&��BЪ�b�l�S�A5?���qZ���>�զ��\>*t��g����AnH`Tǿ�P��gn�ypr�������F:�N��UO�*)D�����l7����Wy􊯻׈�7b�J�VƯ��vA�6��(]����uU���僷\2��G��:�����r�_tn)A��s�X�d�C}��9i�)��)�K�"��ߕ�x��D�La[�=��P��.�yƇ��-��HZ����zپPNd�ˌW|\�V�<w�����r���B���D)�,��*?���\XL?[��u�{��f��a����$���3;mq�A����֝|��EM#ޘCY��5�-��x2_>r�^�t���x!�8q	<�N�݄�+�틬��݆�fo����/H��%/�_��=�ꓸ���k�tmX�oS荣��[d�����kZ9F��J���D��|�r�C�`�ojeS�"Ĺ��/V�UK�)Z��͑�]�sDN5����N��Ɗa��p�����aY�FRzl�ל����ۃ^z^yF��3t�FRvM�$U��<	��DX;->�d��_g�e8ݷ�7��eCEK��u��递|6�i5�h���0�=�H`_�	B��y)VY!��:�wA��ɧ��Ns'�Ā��}&���b̾����/n}
��5���JZv˓EDH�J$�ړ����x�yl�x����;�,y⪩���a��/�m�c7]I�y�|��m��7�v���ɫ>v�뙙r`	e�_�]	e����X{�EL��#3�#�#5������s�v����ۏ���gWi[[�����X�5:
�7�x��=�my|E	�X�U��2w�g޽:Bo\�E�ۏ]�r���s|�x��b�����V���;a6�~��.`@��u�����W����6YY�rBg����K��Δ_I+�,x�U^�����=�v�N����5��b�����I���:�a��P��_n*���ؔr����{c��	�h[_���^�+��t��g���~�Q�_0��VZ}/���'�Ѿ|�xu��A�k�Ys��%�LQ5�f;W e ����|�
V�%
ZM�:��砶��|\�I�	!�&k���t�..����\�+.qz�k�Q�HX��[���C��<'��hp< Lc���-�K+<�ud~���vf{D=6F��ú���>t�%oG��<>����v�	̸+����L3�B���
 ��
��ٯMm�И�M��.�axI��v��:_�6��k�r����IevQp������j�[�}.i���E�U!�q^g�ɯ�^�|eHK�AbD)Wv�U��~�aX��v��ĻBi�˻�Ƿ�6sT����l��ި�$�G�p4b�/��)��mZU��Mζ�Υ���xf��(Ú�����Z��>�	��T|j��i�d��B�����T�%�/�������?����1Ն�;ü�#5N$G[@)f���������9��&[>n��`�'&Z�t$Z)�ߔ�C&�u< N��;��P)��D�i�K`�����&*��	��®�C�H��S�3��-��s�Hq�.�?�n|�lC���:����(�YQ9B�k����ԹMMc?��cş-?�������3��p-�`�����(g-[�م.de�j�S�g�X�9�����E�+nZ:_���[/׬	#{����b����<3v����ţ�1쟡����r:C!Aр}�M'�	:i�O�zQ�Z_����V7�즮h�>��M�=d�Ȗ4t{ũ�ݶ�{K/��u�h�ek�Rb��[��kZc��]���·�eo�v��$��`�$��V6����U�<�)�ޏ�/���o��X�7~����P`AYI׻�y0Գ�H�G���Osz*��2D�ܶ�F��zo����1�0� >2o�^�WO5�}���E#^f���8�L��'�����;:�U.4$a��r��m/�չ�q��o�෨1�o|�R�B" �_�L���CCvg�
�/�=[��Jj=��YD��d�<����ܼ����5�<��憱�#���C��t�>��}B}�^�;����*/3���h޷*N6����ѕ��Roh?t�PFP����"��.��r��K�@��>���;���3�[����K����h}q�A��}�?��,*!�)�ŷ|��$���kys��/�5C9r�iӫ1^�ĝ�t��������6�]��oe8�����s@[��ϻ�=)�U��8Y�~tHQn��B弧;���6�ԭ����RWR�4���m/l���z[x`�Ur�9U�q��G�� �L (��}T%�y�߻~�x}4 ���Y�b��8e�	<���^5�Y4�����ǅ��:D��'�SϢ,j�H����%E��W�O�M�4V�.�.�8��c�94��w$��+��=��ז�B�<ěz��5��QK�4i���P�Ibl�.v<��c��E��c�f˩��ԯ&
E�����	ƿ��Uq�Y��nƑ⎋�͋ �]0]~����u��(b�v���&�9��t�n��%��dp�}9��JJ�܅�4ܹ�n��+���A_�̡��Qٻc�%���A��^��93�x�R����>d�i�3t7�8"���uo� ���FY�/7�f_O��]}n�����y	X��6���������䨋�<���|�O��>���z}xV���+ ��x�z�>��e�f����;���f(�L%���7	��tT`>�YF�r�U;f�2,4�[1P��KC������y���mi�%K���|\]J���R: ���0�ӻZ�$�Ʒb��^bĎ��XO�"�^��H��n5N�_݋��-�P��*ѹ��7�W'�4��O��*zͣR��#2P�X�h<���mm�|x�j�`�%�Y�s
��<T�N�>�ݠG�u���x����W[��	M�~
f�y��Jz�ʭ����mz�����+Q��Cmv�\����j��wM�ɗG-h�3�d�a�-�!��oe<)���Ϗ�g�fkf�8� $w��:�#r��ʡ�C�-؛����#s�/�9U�#i3�����um��uc�]�ε��=��A����OG�i��a�~�{��������(J����z����4+O&�L�����[�Ѡ9�o- {X[���=�6�jO3��W2�L9��c2U�dT����ǋ�]/����K_�c~o���*��(Z0�ǜ�Ė����)�\�=� bW%��(�v�鹣�]{%�|rr����	4�')�ȼu��L4��z��xĤ�������m��O��F���c
����7� ߽98P��H`<<Gy��7��
/���b��A��񡷮��g�>Q�9�d�2yQ}y\������#���C솣x�}=�Ѫ��V8|��N��A4b�-�[�^�����A���\��/g}���^ѳèX�Cy����^��y��m�����`tl���{�M�D�S�.��Sk٣�oW����̡�鹩�Emz���y$�Ǻ�����g���J0!L�R��f׍и��خ�	0�SL���oSO^̬#ђ�+x(a����^�tm�to�d���I@l�g[)��&�_�q��;q�����=�u˯�R�M�:��Ǐ��j�y�S���ճv�	5�w����P<�m����5�mRb�s���������\�t��"���Ǖ�i��8m�z��M��y�y�W� ��-8����V����xCG��^���_|�K���Q�� �y��� ����\�_��ʾJ\����{��6V���zW)|Ȥ4�_����9)`� �:�G��?�K�@L���e9G����ڹ�N�V4�%m�.�P��i��X�D�w��^�e�5�*A�p,�N����A���dIF�y��t߂i`�@����c�3���wW�X3����-�O\o�%ͷm��9�2��?���v;�A�a�1��ߍx�\��?C��+�A��K2�U�����|�(�]R��hJ)G�4��	{s9�ݛ{P=�e��r�6k�ݵLv�Ik�떺��ͽ��p�-�����N7ڛhqυ�OG��W���1����9K�A͆�!*$�(.�]�	z��k�M��;e0J,�q����ўf�Ǐ+�l�%����k�5��6��f=����=�A��ˡ3J���=g3���U�_s�>ُUD���#N���S��u'O�v�h)<�<��݊�04��+@�\_�4Ԩ�B��F~\��^�HhDa|[6�n�^O��X��7��� �f��8`�I�^Z��LYk�1���w�7>�n���;��b+��̃�x��+���\D���,����)-�	ԭv5^��Q����h�%+��}�;]�K1��p��x~kb��]��=�H�]>���ӕ��&���g�~y���?R@��1��0��\h��XM+�	�j[+��b)t��p_z��w��x�|sW�7�W ����$��ң!�,�b�T�|��ٽ��nD�A�R��P>� ����s4X5�;OG
�=�fqڷy7AU+��_��
U�{���ȏ��{��/����q��h��6�ϧ�r�1�i�WiK�G-v�����k3\��?����3}���{q��c:�e,�Y@l�$���x�BOhF�䰼�iU�t�q�}|����.�ĭ�[��v�YNf��^���}"(*���qC=���F���;n��9m�i1�/%�LƄ],ɐ�l�a?��ͪ��{ό'�#6M��w�{�J��n!.8 �$'�܁�h_]��0�S>�2ؾ_O�����oj\E|�R�H�9���h�Rr�q�[��F���7e@�T���^�9=^��ŇS@���(Y���)�#�\pn�خ&��$/���ɶ-el'o�(��L�?�{�w� I����"����aݶ�e6?��N�I�K|�[�^�[#(뽴���7
�xM�	��d��f��q[�n�Y��}l�$�ˏ�M�t��tJ�ɧaxS��-sg���h�iZ��6?��4��?|I��W�R&�Re%_Ѣ���YCQB[O���$����']ǘ+���[� �eQ3Rt�|ڸ�E��$��1��n-�=���=���K�ٹ̕���M_'��&`�Y�%��G�R��跽(GKi6�<����s�С�"���}���ف<�������=��N;С���xNT>����ļ� ��|\Y2�G��o���6��%�̱���v$v���J�}����u��ܫ�����g�����sy��/��H�M[��* B�$_���3�i ])3y��-�����D�W��Ts6�D�9����4O��Cr�M=*tJ�/n5��ٕ���y�c2�s��%��`���>^��[m��*M�9�S����ǲ��۶x?�;�= \��G%� ~K����+�A�h-��tu�e��ǙCtӕ7����� ږ����Lď������(~?t�<�`�C%A��S��R��
�b�!T7�H��8[b}"u{g� �d�>T-6|��^}�&m�]x��hŹ nAG��l+vR�*�,�[�c����R�h�0�6ĭ����Ȏc��q�#��R�8���w��!+R��חۘ���1�{�}��d����x8���F���䑩
��ʖ�<&�Wh�������d��Z�ksS�C����rC/ǫ��G5�9d��`���՛d^����N�����u�?�v���z.�%[�����s&�R�ΟEDl�T;�P�}�D�]�*1 H��)��֢g�¡d^D����+=}g�-7���*�-�N0&I����|�ې�+ʴO��n8c����Gw���
_<���Gg�d�mq��-��>�U��F_���X1����}KI�s�f#�z�����)�D2|$)iRW���Јd��'aMaG���}}|S]�^M�Km�+:���U��'�3�&�j��{�E���_Ty�� �[Dǭ��7�n3]�ψ���r�^f��v��yoQ׎^�g���	��J��'Z���\+������^�����3?�_I�r��
�V<�����ϗZr��[���e#:AG�������=�����=_�c���]p3r[!筮�V,�ǫ��q �M`\%]8+SR#U����i� ��I�s�N�
��*�%1�CV���A�s���͖r[�Ƕ/��Xz�#@��p�x�	T����Ķ�J�dz7������ݺ�	5-9��P��%��=�)��Ϸ�	U�s#�j���}[2�w��e�g?�9w��y��������/�a3�}��R��?z 1�ⲙ��
�;�o�Lvm�DP�������y՝��f8�������R�OF�b��d��N�k���M �R�h�O��G�(��{0_nK1��ʃc��]'�:ˎ�4֋O��<�ߜP�$[�_�Ik	���)�9/�
��������O��q���x��o �KN�'e4&,[w�GbVl �TY*�u��5cF�����m���ݚ����i����ȐЩ��w&E�Gh{������v�o��'��3IRG�}T��-���<��eoi�a�XH8�8���1|���$W�dP�)�cO��I�/�����v�W)����]tH�IeU�/���~ ���#=w.���wQ�[�?:3�<l�br�� }����ʥ'�)�&�&6%%�b6����5��4/�~>�5�ݷ}nZo�Ж�V�6�N9F0E!��~�6D�|�}YG�`HX�&D���$��\<��<3DQ��U�jC�I���ړ3o>�����
%~߿��Zc�$��@��	�l�ϫ�IM�d9�y��;���	�I���:��;�ՇI����W�~����ݞY�6�W�
��j2E�/~^�A�%�#?`G[������
��O�P6>�ʐ ��Hp6l76��,^hR�u7�
��������;���Lω�~���.s�"ɓV�_�1BHP�z��ȹ]����v��)Ĥ�����E�\0r��;.oW�m�˒�b嬜�΅MA���\�;�����&��������(�W�2U@�ƿE_��j)U�-A��P��'��d���T$�����9v�c�M��N��拀ϯ�z��pk���I
���	&hI�(��Ӣ&)Xx��ă$@�.>K���Ks��]fY�A��j:�c���?�ژ%=d΃�'YKm�u�^Ȇ��`R�D�zB�ϿuB�Q�;0B�gzTa�ku∀��n��k�>f�F!��=�D�㟘P�>��&R��հ��cmLwT�od҃����o�k:9D�N��@_�����o�Ko�r�r�h��ڔ�D�-AP�M�����Z�R����)3�'Mw\i�*����7Ω�������^���l	}��.��.F|�͊kϛs]� b�g%}�6��㕟[��2l]R���+2�t���Za�s_��P#B�c�}v]�mqFAyV_�e>��H����G�ѕ��¡ɋ���Lo����h�u���J=�_�b;�~)Lt��F��/�-��URǕ���̯�s�)G�����7�D�qN�֗��]����4�R�峴�����o���׏�s2�x�#�	p�,>ЙF��2��z�h�zc�Y#�	�8)7-���^e�o+b����˃0M�'Ԏ�s���|��.��wŰ���X}Hv���	Pe�j��%/ⷬ��"�9=!��c��ǃ�>�C�/��4��[Ⱦ;����T^���C�����DXYL%��u�^��^l���P�����̻§j��zIXH��j��Wp��@��Uv����ѫ>�$=L�k7�2�vH]�
Vɟ��ξ�:i����e�7��8���;:�n젪��c4D�E��A��>\����[��>�51,�Kd��B���g�TM?�S���<��O�����?Ő�3p�D�C�Տ����6D{T�B�-]�vLa�ј��ɺ�%x�'q#5��+��)d�����\�<�_Y��� �_�>��s�����e5V/lP�y���)��ԫ��G�8�y�)��r�b��9@x���Y�c��I��97�_�����|Y\��|�!z��szW���O��;�<+�Vie������z�@�fQ��U/����1W���v�Aw��q�H�1�}�����@ d4������EUՈ�*ŷ{ceT���X�aRt1��_]NI^����>��ݡ�խ�Rqt�}�W��a�q����sV�}�C�K��=�/�����ruoƪ����yS�h�E��u�<�cr����-|�dcت�k�Ա K��/,8�\�&Hi��ō�ٴ
mN�+��k����m�6e=0���@����R�l[Z�Td���Z��q�U��*(($�Z������IWF:�Y U�tP�YW��9�* �y[�����.�*�ѩv�CJȏ�*8ƕ��r���� �7���Ȫ!�U{s��M" �G���U;�;�(���w�eTT�
j��\��)U6A�#V�4�=��w5�_��9Z��v�����_Qe�\Tk�*�*c�y`���
B��\��U}� x�_�ve��@�N֗���:+UCҁ-�
>�����K�0����Ou��ϙ����>'�P ֩���#[�J��˧8f�-��)p8��}��B�ճ����mv�j��\W���!"ۯ����kL�H�|��>}v�M�v �I�̽{�._��b�K��	)CS^Ap���\���ҌO�B`���a�c,jwr)�Ҡ����>u��t�٦� S��h3�~o����0����X�����UT�2��DR3[��'U�R�tᩗ��D�2E����H�����V�@�vXG�J�����ƥ�lc(�����⾒��-�X!��cJ�ms4GO;������Ƀ��� m���>>���@T ��R��d�CB�$�14y��������I��t���#�Kc����2��|����!�Y;��_�]��\��(�X5�lP�t�	rE�|a��A�Y˒&�ɝN��T�B��4�/1���rۤh�K����|��(�M_-��E���#`��S�x�]�x��?�v�>��9<��PdjH�_�=�A�-{>��f�F=*9˜*""j��$�i�j��xu���}�cy�zs,�	=)i� R�7����>:��ASk_�~e����v����c�(@k����b�Yy� �cP0��z�����{��*Y��jY�Ri[�x��έ��%Uݘ�
�Qօm7�G�H�����v�ܵwdg1+5�y���\����]���H��3X��1��?3�b�(���x2_i6�CR}�P�0���v��)��e{U^df�ҝ]����t�\�*sa
E�Sj�� ��<�|yEҹ` |�Ɗ"A������$@���ӈ�o2ڻ�i���%��Wq�o���/@���w�,b;�r-rB�.*��J�T%'�M�����'�k�?���73]�^�����T���c@p�F��t}�E�%%:�KM�s��1�e@�Qg�>����ҥw�J�q0���
_W�����ƹB-1�[��˃&�}�l�@L�ھ>��sTul���-kFLQQ�|F�Q�Ӆ}�!�g�i�1M�ל��mb]�~pv8 ���Wz���)���´度�Vi�.�hO1ɇ*�lWe���\$�ÑL����稔�ȣA� �Hd�-�,՟s��F� ��A�%�2+{�~"$8Q��!��wy���M>�w���5��o�#�� �6$�����r>К�
i��
�[��w��P��&j���5�r�G�8��tY��.��bQ��p���瘌�,��_��^�n
��;�x��C�-MY�c��<c�ܼ�&{���S�s5������5t'���H�����@ϔA�+������l�{�552S �W�M�ZRTЉ�oEy�:�л5W!������Tb�	V>�nϡ�Zo�{�p��;/�=�Oׯ�T����xq^+�Ų��]*h���P�����[�����H������j�����mmA��S˵�3r�%�K���][kS�3��Bm����'}���;n��ɗ��
��%�:9���B﵅�DCx� @�j��Z�VM��w�H�^#^ ���r. ���R M5+W��ӊ����X��|�w7ї +t��jȳ���>�d�9�C����H���VxQ���h<{v�k�L�)��v������qC�h8����UۄE���!���ǯ6qoK�̦��Y+Wgޑ�[S�:�LE��Nu��(n����'�����x��j��\=D5�~��A�G��Q)WA��ث�|d�� ��I�����<�o�;�9/�َ��S�u�t�{߃�m��>}�ԣk_�ii���o�1^��#�����X��b=���&l����S�<��ǧk�"EU.��qM��SL��<5B��p�zL�ҕ U4�y�#(˴#R#[��p ���c�y�G ����ְ�p}�FiJ��l���������)��0�N!��>Y=�X#�`D�{�f%�޵��&��T��J,z�-Ȫ��.c�Ȃa@9B��C�@���%1�g@!� ���6虒��tD��2�Z�5��R��BϟM�����\�X�_����Xd��NmZ5$�^�7Z-Ռ�|����ɶ��u��򼩩�ny�q/���ǃ A�|�)�V<0D�4⏾�_(!��ڣ���e5����!N�|Ѯ}K�rS�`�If �)(�ڟ)���� �!��y??+��:�a���<V��ګTS��|u�m��𶴲��{\��᢬P�g�!e;D�y��
';�������N�a%�w5��O�����X�Ţ^QQQ!���� ��h�AAW��C~t���T
 ЄD�N�Gյ������ �wD�d�dgg��>}�v �]g��.����s]�ԏ��I<�u�( �xZb�􅈂�E6�kS��.����ɹiY�I3���/�_�'�#��NE�BI�����7\����jJ�&F� ���?��\��?+�\+���~k5Z�"�D���7iZ�E[|�?/XV��g��$�L��k֗�\����j�Ѕ�S��}�t:w����?b΃+N(�������,!�O�@��H��H��wH�k�H3A'Al<~�b��Dv�t��v&�/ѣ��5��Ը�j�7(���'zٙ/@=�x�n0��ϯFKHR3#l�T���
�y9�m׮ ?�HqW{q�3Zvg�C�tXWVVFt��{�����������7Y�k#}�bc�?<�e�1Mf�''Q�ش>m�b��"��ᡡ�2���r0���D����?���J�F�Q֦1\$}���24dD�L�
M��F�ɂh��ɡ�/�B�6}�;���շD,�e��kp7�5�	����<�xc�;Dm=|ҵj���`�po��ؔX�M�f�)rx��m�`f!�5������ny��T�%>קaH�a��%�OҜ�4+�{d~��2���L}��E�S5��� �X@�$(:�;�K����W���Vw2���2�]��ܿ0(	����`B��[FRQ붳T�څƯ�V��M�=)���)�g�;	)���s�R#y�݉t�cEF��1ve�T__��(����¡\�x�d�0��y�o�2���B�H_����K����;J:Ƌ��#�!�_��*L�$��ē6@ۢ��(y&�5K�I�q8Z>��|�#$,=ճ���.+��qL,,�t�B6��|�J1��+���\��}6�9�mӝ]�����Y��W8b��b�%�$d�`�%ڋ�wc_�:������C�>�ݮw��q���m��I~�lg!m�6�-3��В�e	W.���(��� �؁D{F��D{���l��Ɏq ��%��<������V�o��?�wT�8�פ����(�#b3�Oxt���Ǩ�����w����V�����cS83Q;j:�>_��{(���8�Hh��E�����ǘ2�5�7�����?E	"��x��S�H�"@�F$8Y���|q ��L�v���=@ �n��v9�1�N�F��dM����w���{���u�0�
�Ҳ�
j��;���P�� �sD�
�**C1�W���%�W.U8��a=�Y���8)�ç����	��\\�D�+J1�t-,2����2q�?��f�Y���9�/n՗N������Kh�H����߸C"'�Z%:�����%��ג�|��$B|�!�T=����\ jF J�kl�;�nuH�@J�1�ں5(nN���z2�4��dY�������OJ .2\��i���}��&���8�Ǐ���G����;L�H��Qk��1�A�5��_B��/��Z�u6Y"l{Ox�S�&A]�ծ�E5����C&q�gV���B|XRؿ�<�+�n���M�2�i
\�0�>KY�q2T���z\�g�fm��������Yi�5 |� 9(�,%F�+W�.�����������.�ضv}է��U�W������=w�k��a���"����iQ�����:|���T�2
V|�L5�6���i�E7<������#:>�g+����![r�ɳ��>6ă*2l<;�z?� &$�� ʛ�N�9W�|�wǢG�l����S�1��X�������ؽ����R榰�
p_K�%=?�M��1<Q�:r~s�c��↹0&�1����%��XMT�Ηr)F�G��`\��9��a�9���v��׳^���j���661Ϳ���=��QX�.���g��&���|�o����-�*��o+	Y���>�f��5>PL�/��i��
�|�e��.n?���`���Ms���g���_���f�����H:�K|��Y�)�Hn�笹}:E_�e_�N�����W�C玩.��5�7l�_r����$�g�mCQ�ޱ"�ι6e����gRHR�Zw�G�e�0����WP�VD_�5���L(������-CYz��38�}����]�s���N4���P�w���|au��Ǐ���Gk�|�
>�f�`2b(�4lk��~��p3�U�gKԱ)�;^\w2���(���I��_�������&�X�Y��d͵�V#�9;^��E9�F42�̄%���Z�+�/�9�KD��=n��0S�eՐc�98��bvS�g��.���3�&)U	�� ���)4+�4RMl``�ғ&�f�;�H����8���!�i�����B���E�,���y�}���y�6,��ųp��<[�H�-͵�ʾ��K��,vĐp�q�b�0Zn�k��p��=�5�w���!BO �d��fF���Pj5p=
	>JX�Ж]�ƊP2���i�E�rs���� ��$�4�ÅR��,���te�Z�@N�E=�}�6�e�ࡋ�FD�5�ܹ��0T��R�7�&J�2�m8�|��m�s[����
G�{Zi4��j�E^4��S744L�	C��n�fj��WL���\~�Ր��Oh2��@v ������[nWI	_�6�x��ּ�&0��Y�)��'�%>�t�Cm&R^;��a��~_{�DHL�#��}G(���ľg��	���ZL�d�l�+c���d�	i�,��W���g ��Y�/�2���ԗ�_���8ޑ��0ś�C丂��YzYCG.~~����\-�*$HD����Hq�^ � \bd� ��D��EL�qq��<�X ��x��	�`�i`��Ps�B�݌3����_A����!·C�i���ie��K&M��Y+F�$�1LYL�OnPP\)k��KG'�\j�J���R!��v�'fk�r���������8�4m����eVE�^ջlU���7"N��]|���}�Qc��"W�zpYtu(?ߙ��9�!�Jۈ Е�>P���#K|�D�ԒE�#}a��k��45G��`�A�F�����N�xS��k��[J�ٜ/�י�y��8���,�Y��G?bG*_��=��&>{V�1:��S���HG������djc�k�@��u3��եO#o�ҤW���.��~33���n�G��?�a��p����u�G�Qc�� jgA��$*�s?^5�Y����Z.2ͻ*)�K��ƹ ɗ��eQ {>�K�׆g��ֿ??�GH��/^��D��T _�2���ױ�q#��'=1p�$4@�
n}}��P��=��`��a��aF�(~�j�~���q��
>[�vݞXOSn5�N��=-+ݣ����ȺMMh�T��j�����^�"�>��|v�����$�oc��Ç�r��O����	�J�_`���Kz5��hSX��ŝED���d�"������Jry0u���&����b��Y��.ko��R��/��n��+r[#�r$!��;KDT��zD�|��*��I¬���#��a{ؙK��cb��^1��v��u�T	E��_� ��y' �[~�������%��=j���r\sJ��e}W��I�Ӊ�xB�
�b='���8�3�7É��}���N�7�{��עn̹��:���jAT,
N��.�T�N+3��Np#�N�a�hВ�R7�@��� ��I[�sJ�"��Y�A��"J�z>	���e��ྐྵ�g�2�ۯ���K�V���Ԃ�C�9i�[�*�}��Ar!n*r�A�,/��"�C�U-{;=�������մ��ܻ�M"�~�񺻏%��
�V��j����]7�m�ט�|�#�7�ѣ�����zZ�C�U�z~�Pk �z\ ���~����&����;v��	�j�ޡ�\&cOZcp�Q��G��omq_���Z���)1�He��Ɋ��Li䘏#\�iN���gpΫs�K����=�ob .���F+���iw5���u������E�ls�کz8������M��q����㶧�^�'{����5[Ēǻ}t�������,��ݟ�B=��Ѓs����~�����=����n-o�'�5@z	Q$/Rj�Z���ݗՌ�-+j����Z�#��E0;�ǯ�8�8X�k���ͷ���s~`���`g�O>�i!���t�Ld#\h��� :���g[eZ�Ӭ�d�q'_������p8|���h�|ߥFH��	΍���x�����hD���FlHHH�QS`o���󡢋��k���&���~ӕ��=^���E�����|�v{�i�BhG��v_v�r��̢���Py&`a�Z�w4���~}��h���-C+?{'G�u9��g�����$������kh��%>��Q:|��7k��$�^��� C�[�n���jݫN+��$ �5N�.�j˙�߳ԛb�������v�W\BO����S��ɮ  ���԰�����N��[(�/ �[!�w|������_`{���M��r��b�G*KK������4=���p�1,G���nwު�D���>��Q/.##�ߔ�[�w�+��.O��|ΜK$��6vB�j�b�
���=b���r���,+��4��M�?Ca�8���h'9�u��Ap���_{%d�+akl��]K���PP M�屐�z{����>����[y�T�,��(a�����q�������8��)�0���(��T�yj���x>�h>:"�k>�.�5x=��f����S�C��7 A��F�I5Z�#Ƒ�Ѵ@��9PT�'������[=f�3���b8"��&��	k���l�,��F�,6x��1���|T}��}���Y99�*�V[���F5W0���c�݁���4��̂w�di�n=Y��59l�\q�j�:Ͻ�����
�A�L�L@�#�H�X�`՚��$5��7��qp+��@���?��rrr;��TN���A ۋڔ��̝#��[o8�?2
��%���wZH���jd+�'v�;L(���K��*?	������Uy��YrՉx~�&�dK|g�4��n1��y�m�P0����u�1�(�Uo�U2��up0�χ�s�{�G�(�h_�U���;cBٞ�) ;7[�|ݗ���ʔ�~0���u����W
�E�� ���N�$�= G�1��i@8$:ܕ.��^�r��:/��V�(>�z�ݷ��	ʥ�<����������s�l����8?XL�o�����;�E��19��t�����&�m5�p֢��!خ�T]Q����͇/���<��yR7�-r�G�6V�ٛ�!+V���J��JJ�ۑ�!�y�Ȭ�-�F v���2H��t{W���RK>��>�7� ��]IT�����A�;�pbE{�A��C���kd��D=����^�7.�~>����`������1�Y�����K��yS"�婢F�KRP p��m��>����;ٿl����T�y�Zf���"�Qw+Row�"�*�'�cp�"@.��J������i���V
U)�4��%���goq�Y}��g��b��_K�$ʡ"��犆�WU���#��)�?lL�+{���i?Qr4U,��|B��n��	^�xe��_l
��S@o�H� :���f9��M�D<�8�!�$5�%%�2ہZ���FF�oĢW^Y�%���y�(�x?�|�[1��u!� �I�|��ˤ���5�z)9ɣ}�t}£>T�I@O	C�ek��������V��Zf��F�0#��!��@k�HEQD�Ϫ�߰�!��c�c��}��3)1��H!
"���0��AI� ���H� Rb�"!� ����tw�t=�0��|���|���D��}v�����9�}k�>�{f�}1x��L�y3��]�W8Hr�w%<%I�u���ş�<�\�^�M�ܞ�`1��G�ɇ�-]r�-#(4s��؋��h�!�+l5��/k�OG)�y�;:��Y���Z���!FYeeQ{�*��ɩ�޻}�q��Aq�M��L�W��f�F�ISW�~p^V34L,8G
������h<Ay~�1�*���m��Kq�(MN�
p3"f#�eY�;*�������l�vk��ˍ[��U��Hv�P0�*�O�Ư~��uy|zG�P���F3m/�����f9�<�'��/�"�٨F�8څD}�D������R��@�[.l�AD��u��ʌkV9���՝_ۓ�y5[�Ҩ�� S��	I��S������桸�J�)�}��5����B�6F�?���2Z�*sRIFm53&V�*���V�IW.�����(�Ǆ����P���z鋱�R����(%u��p��8@�^8E�?��ti�k�T�[�0�W�Bb�F"�R.+g"_��w;�f��XTO4��YB�/&(^�<��q�#��G����?~�e����չ=7B3~��t�	�6�	�>�i���8�ؽ���{+|Q�1
Ԩzl�ύ
�$\�9���֬ᐈ��|[G��@M9�4�!�#� m#�BKw_�F��H�
����r�Ӌ_b_�e��e4�J���[j�8Ze?*2�V�pL�04��W���idE�mN���y���n��m�g�������*����y�-Lа+�E~6t�Y��R�H�q�U��o���c����Y�1���#�;w�y8:)��ο�L8~��[<���i�l>���Ю۳���#�G)�Ч�X�5�s��SM&�������Nǈ�.P�� ���%�׃�+�t���ߤ���R�`�pB~�8Z�O�H��Y�Ό(��(��@/��q�}�Y��=�����G?M��EBE.Mmm�[����y/��l�KNo�HMn��-�eK���h�~��F�V�ş��V���y�!o4����㼚��O
��?���-g}���M,��L0�X���K ] ��,���MBdE#�	��H��̆mU����P�c±|����sJj��B�'�0/{���d�pY$��󌹺��[�5P��";�j�����k]�>��z_����M���Z���7��A�#L��\���Z���+�����5D� ��`�+�t�,���Vx�# ��Mg��n�l�/<ג+�C�}ӶIv�F/�Ä(X����4���)ϔQ�e��}���˗4\����U�i �̚Ż/�,ƻ��[vs㟎KR0�儚2��!H��Q��H�r[���!���zd����sWlw��ϛ��ʦ^�}G33��� rQ��]��/�J��w�Ѓ�V�k���7��o�z�lq�_�2;�� �OV���M&������T <d���M7��iܥ�Qγl���'��5q�V�zr&�^���
��FZV�G.b;����4����l�u�ȎI��Ω�C���ᑷf�:����u�4�a�����o�Ez=QD"���~(�k������
�$UՕ4�$kjdD�ȃf��]� j����/"`��G5R�u����7w�`i��{���]E>M����m3n����1acjn��Y���ΰh��6�f7^ACJ�Z۝�W�U�:��S+���gш��u99߂7��@�S��d
�l#��f@�o5�>����8(!4��^�h��#�& ?/s�ӥhg���)W9�8	�*9XKn���/�sq�>�m���#��G�.��}�%�f �w�i��J�����[2�|���Օ7&��!t���PO=�t~�8�����c�u�6x�\n?)�M�zU�8Y�]��573���ڛ��b~���������Kp�/fw�_�acɴ�%Cyw�q���,��r^������H�|A	Q"�4�7��`ɐf��Z[gƱ��ܳ&����~��Ss�1��D�q �`q>Nv�}<�k2���k�K�d�����(�,N����P�Lt���P@*�S
�Ҍ���ßx�V��`9/.��@�����NBA��ZU_��[��L����M����)5կ�ÏLw�Z�z&�,Y&ǐMl��6��ÄQ8J��u�r2ء��)B��!a��r��Kh**�	Ɣk�؞�B{ňXe�8,���_����ܟ�d�Wl4��~k��S�(؋�@q�]�s���v���>R�X%I���#oK���������i��D�q3��wnc~3m ӓ�'�^�T֑������nn)z��Ռ��
���'v�I�I�=�{*ֳ��9��Ok�8���D~5 �}���x�S
[��~.�V�"�Ö-AJ���n��|��mP{�X3��g�����f��M$�pp��s��XnIe}���-��d� �Xr�92��,E�D#ihE�� ��Vn���|f��h�%���UX�c`�z����(!NI�/;N������:=���DĖ��uHΟ�@j��:w��)ֵ�p�I�����0^z'{��՗�ϩ����u_�ׇ���;A-a���%Z�۠?�#qg�4�:�+'8�5��m�%G�b�W����!l��Ŷ2Lj�G�r�}cp��P��{�Q�b@>�y���9��v[���B�����{J:�89��4��0�}�N���h���k�h��pf�\��w�zD��y�:�.ǎ���Eԧ��\� +��m��<���e2�4^��ٴ�A�=f�	����w�m��B��&2	��4��QbF�:�[���w��9N$�G�	<��ARIQ)� ��^(|타!+�_�ڹ(	0�rhR����Zź�f�y_��Βl�^�We崨�Kk���l�v?z��}ͯZ�S�g��y��пg޵L����L-.fۑ���M�J��r���jڨ|�X)!_���Fq�1KXS�Q�,º��)����Ge=�C��_���t澗���-�2V�R �3E1�1��ϡ)
b�Wr�c�����
�i�?�	Aߌ�~4�yB`�n�R�mW����3�\K���b�_���}S���)f�V���q�"A'=9���#=2��
����@o��$(��L��Ʈ���~ҭ/�<ww��FG����so>�f�6+E�pS?��;I��R��F�׏8���y7�1��M��	<����N814�����J�rvۆ�����W[Yn۟��jbo�R0U�Ɉ�
����Ρ<%r̢��b�"�<y����˗�=�Wӿ�4���Uh�ob�rٚ��R�q�����}˜��6�	�t�U��ڶ�F�,_a!�X4����bL�^)nxyOƃ�Þ�"^���=7���Cv\� �\~.?b7#���x5/oRc�ʭ�yJ����6u�}�v��9���Fsk�B��ͽ��j�+�K�m;B+�z���Y6�]�NUs!0��]�<�qȓ����<��I}��b�p�/d�_��Y<eй��W��8�j��i��K��u�O7��>�0j�oʓ+n�~�����߽GyK����/�B_���.nJh����Ta9���G�P� a�A¬��enN�����o�(677w?V�GsX4d=BM���o�S���[���X�rb�}�p�ö~��M'4�+��Ÿjd�\p�c���}���6�-%�?\�և������7-��I�X4�T�I#�/_�~	A�����=�(D����|�,$E���]Al<�����N�i��έ�ƤGi�kl�'����9E��޹ل,����s3�6�� k�[�֬j�dacs�@{P��[�����t���û�ڙh7�'�l�b>ɥ�+/���Yj�:d���?Mx�q1�۳g(��1���k��/j�y@J��3��8� h��լ! #��v�n�I���ec[��v3�L�pXr}��Xt�D�	����]Q�p�_SI�nD�௕k�9,5�__����ͯ��d<�O�~�|2\�9VzHˆ���N��n��`��4:�-y[��m�&�(nc�4��騄�<on��Y��&4�m���y��pz�e�$�۷���KD776��su�:��d8F�$(-=�ֺ�RK'Vdt��k��Dq^_��'�0�����RM(79(q��Ά�m-�.6�H�5``,�E���� �2��|�p��O��''}r�	n��_����r_n�ʦ�~���~�eJ�奞��]��Lu�斖���i�P�b��(`�sl�����t	l�����:9B�Σ��X0A�	�>A�%_��;m}��\B"��� �0���1������1�	
nߞ2��Ҹ�o<�P�~T�'�"��h��{{6��l*�`-/T�q�����'����.��6��嗌�?7L:CxF��X�H�?"*��ET%�2z�w���&�L+��P�Q���%| 2��i��AQb)aG�.�4���pǞ�� Z]��r"��1V���E�2s�Wшd�?�O��3����f���7��Fu`F�=��J/�$�
س�y�&�OT;�?C�]��ڌ'���;�~#{������s�'�6�b���XS���%fq�d�b�!����,�1q��.��+�Ÿm	����8�~����؛��`͊�7��%�"=�K�]�������%?_�s���w��炧�Q k���W����>#����
��T�c�p��B�8���/$X{�o?�+Ĝ���!��Ē O�o�	��?�I�VyH�##��nJ�(<q�o�y�!q
/�O~��_�[���MAS�>o{�3��D�-�`�r�V�6����4�7�'nx��[��.0�����_��M| =�[��(mY?�k�(��$7���|/B�j�(�<cD��aHd�hl����;A��>s=tN��w١ˢ�������L�1��j��G��c���15�i{H�I�fǙn�����B��7
6"�Щ��ؕ����w/j�8>��4�a�{n�^;�+{���^����S��d˘���-�LS��W��jtj}z����Gj4�!��gN���U,�P�h��끁�#����,����-`w(e)|w�1-��&s�K�T�^��>�/U'�8���o��U �fax�}�\<�`���p�F��z��92�����m)Jj��)���)�^��	N6�A��zh�ĸJ�\��3~�ß�U�ylӿ�a:�4�N!a�Jd[�P+�}*������b=_�A2�\�Gr�Oe1DD����wB�*����� �����^�J~����1SԼ��J����U���L�7�5�S�~�����eq_��>�iw�,��2/�ϟ��� ��2~A����ʵK��Y����(��|��K�s-JEO��
\�����L��~o�[e�륰�����Ģ]l���i�nZ�?�6S7�|`�
���4��:����(Ő!�ݧ��\������6��߁��8��Bl�f�IЂF��@�dH��;����f�Ը�Ƭ��V�x!��v&'7wvh�3��6�^����m�^�d_� ��3YǼr����%�Ȉn�����s���Z��į��[���p�IJ�װ *`�Z{x1��/�HC�f�������?z������m1�~4�8��
<�����@ܞ��B��ƺ�^2��ѷAEs������7��QoG�	�I���>�d��)j3���*	Rq��33�K�D�Q�>����!'�+�S��]16�[�u���O@��h�i3���T-�%:Nx!n���*�YŌ��S���=x���_��o��G���sw~{�����>`dG���]���_�R��x�z
S|xyJ[!R=T��-�<�~>�F3�s��Q2h��T�r����f�v	Y��8|\T���b웸�ccg���͐������}�3N����g�����$�3������r����	�L��J�m����W?>�@d)>'h)�u��I'��.�oeh(ЏJf}��p�<�� 8��B���b�
K���H�"+�?o�,͆S�� m�~��o�k�޿�3*^�~}[eǜ�;���_t*�aM�s��^�����,�����U�5�W��/7���Ko�p��&���ō\��У2t� �f��n�^�{!��]�-���'5n�/k���kj�K�������S����R�{!�#�ڬ0�o�UlzD�P�4�&����`�l��auT�k��d}=��i�"Z%=��Qہޘ�Da�a��g�ڞ4?t���b��{z���R���1O0F��gW����ܻ>�=��ш�~�t!�]s�M����8�����G�A�}o��R���L�bRZ��c�?f�F���<|��m��0E�ܜ��w��˩�=�Fl %��.
ըHɬ�AӍ=����m�X%_�H�Nˡ�����������▊l�tSb9$+%%��qGۃ0俻�B�./O���mF�Z�~������4�ϴ�OT�<�B�Q�mP=�0��O4	��<Zޯl��rf�J!����?H%���~�/D������o�܋��_��e���	!z�`T�5�j5R��gè�l�v���XDD�{<�#c%r3���+�o}����mĻ+Ƴ3��r�͉���{�7����bv�'|�&�Wt��r͜An���<�8񢰹Zq�p/X�?[(P��r./��r̻�����.C��1ۋl�9v�jd;fQ��=)��?�-7���;m������uƧ��h6�H�I�y�<i�ki����.����jx��G��Z����T��U�x���>H:����	�j{e�v��e��Ňw�L�b��!Dg���������H_��?k��Z��j�ְ�v�h�8H�N����ρNq��e���<�Ҍ�*��4�/]�q�COQ�'������I���#�%_�3��=�Lz��\�o�6������)��΢��
� ������IF7���E�󬟛uv�&G�����_D	lA���S�{��?0�����d:�	%>�"�"��pDO�K^+�u�y�c}�)��R����'�������u�s��2%��5�NSqU��>��O"h��,�܎t]u�>��I�`s��LMG�R�ʧ+�ם�Y��:�1���w��ݎJxG�od�o����9d��_�*wE芧��Z�6T��i
�>n_r�� Vb��
����(чC�Ŋ,��nM�O�Fb��r���y�\$$�V"��v��A�p��@�YZ�O��� R�Q�P�u��L�GxO';::�<ĳ���{�ꉈb�K�X�����+�L�����/�h0�B_�G�%��F�{��@ �d�i���ǃ_�W��\VO�������o�Z�'��
���.30^��-�9;[��B�R:#���'EOx-��W�Ŧ�� ��W`KK(��M�����~�Q�� y�+E��}[^�Jc�#�2kmW�툮%_u�af})�/�!2	��r�ч	Ų����ӯ	*!;b�L,�SG����6��]�-�} �$�������pv��ĐP�K���NC?�^�@�`p>��k�(o��fF%�2>>�W��/�O��C�ӟJ�%�P�+aJ�l��+Z�����\�*��6�+b�?����;�-�8��|��F/�+#��4�^03�e���j(/��ړ���I�����;��S��JO����"fS��
K�+-�{��|=vb�\�f�+����"�v��1�$�.�	���5U*���YȎA��j�����7�e+|��X����I�@���6�=��׻�ggʞu5-�-�'W,8�n�P,�I8�7ߘl�-�"ד�ԽoU_hw�u���ޙx~*�+�}ǋ�r�>�qF�=��͞ohS@��g���/�0ǳ���Ӊ��_jI����+X�����V����M��8$�7�쳶���f�9��h
�EĒ�Q#���^o��Y��R���mGΣ�E�xn���T������Vnp�VE���j�Șō�!���kN?%�"$T_�/�q�-$k_s�wx�{ē_)�.��a�A��@��X��O��B�Щ����M�=�|VQ�f��:������g%��K?l�X&�8�O�U�^�Y���Ý*��\Enʕ���G����@x]�>�3�ӷ���pW���#���T��և���lF��Ŝ�^=ng�fm	4L��]�rV��$f}��=6��,w�K�����h�[�J���O�kL����s�T�l�Z��Mh��f2K�[M�� J���$B�*��p�R�5�2���Z�X�(/A�U���Ϲ�'L��x�p�[�
����Q�XL��o�;m��%*?0DX{7>B�w[k�h���g}�����i�'l���v�
*�Jw~|�����Q�]G�΁�ڥa�9�GvQ��]4aZ3柂jx��?�Y��dP��D��U�#������x��D� �A��&Hц鴋s���a�:-���:i9��T�ų`��j3x-���p�� 	�����n�>����[�j���,8�H���/T��{xa��W��8�Y1�_Xì�k�w�����gØ����	�v/1.b��\o���@�ܼ��yx­0ЅU6�r�&O�`t�Z�d��2�ź���,�:��߫��n?��ʵ���B��G��Y�  CTQD bP�����%֖�`�֟1k�`
�cPfaVF�����- �:�s}����>Z�5��Fy�	F:�r����X�{D��-e)�W���f�E�zf�����l�GS�^h.�x�.[N�ۓvHh=��V'��Wd��v��^7�䤟z��cE�A����_B��;���l�}!ĉa.���5�uu.�Q�ի|a���u�R���i�C�}����4ŉ�=y��>�����S� 0���P���tFe�a��_Uk�|�?Q־���_5C���Wk�ԭ~֡�LȠ�J�fDE]��!�n�� �� �
���I{���n�靨*	J7�s��ܷ��E�%�r�k�o��� b��q"��7�\n��ﲇ���o�[>��㪀�B(�������"ڴ�%�(�9��p�Ih��4���-��[~q\��\mt� y�S��<�k����W��GJo����㱚L*��^� �J�,�\�X�!S#.@&�J���,a�R>Z���8�����Uܳ�\�N}���X�+j�'��Тmj�:��fR�8��_?���|;7ߒM�_����4�P�zP�ۑ+9w��MK�ݯ�@��B<.�A?��"An�	�@�jH��^[��y���A���!s��3��d�퓱H�ş������]�Ǿ��yҽѕ�����&�5]�>�����r[0\s����\���~C�X�'qLW��$L^��t�O�Cc�/�����KƉ{�~��#$!ѥ�!Rvk�?	ۆn��h���y'�<(�/Z^^Wj���I�#�n �}O�?���<���:�U��88�{�&AR�t��Ŕ���k����'���9-�W �BL��![p�i�Iآ�ݡaM����lKw���H�����c>��&�k;Bx���*�o
����C5u�u���Vo*߽s{��u�d˽VQI_Gϼ� Q�z�ˢ��F�m���b��,��V���<}���˙�h#K4��P��,���@�^$�GI<�qg����-�4C8��{m'���~��p�lt�|EI��_��>QL`���-��g�-�(�:h{�(!\��_*|�!������RL�J�x�����kL��s���T0,�q��N�p�V�7�u��yp;_��k�FФ�ݓ�?9�'��nC�EEį�����*k�2U�Bz��fk�����/��N%�ZR֜P���`��[J��A�4S��s����~0��l�6@���B�9���zl8J��[�I�@و̽`����������m��q�;�3�ۏ�u�hҤ�8�z��۾�}]"y��$�Y%ӌ���p�B��CMٻ�C~��^�8���������1��B�pg~Se�O$%��ޯ/|�v�4S�DF��7(=����3���l?�6N����m/t�r�����_�x��N�J�|e񆥏�>^���ڗ�O���h#UiT]��`�)U��v��իq�f�S��ï�P�n
l�R�=�b��r�w�`�`�Z�#��
 ��g�ޢ��Tm6��h68�qӄ�J�Y����{���fk�f�I��Y��.ϳ �K�L~���/yW$+��L�
N��k��ެ�ϝ��t�6��^���/�{��GQ�Z�&�}�� L��tK�ꃱu�����,i\�uI5Z9Ha[����p����egN\yA�f��J��[
���~�F���qO)��Ӎ�'�qwY��n){F�j�b�[U�Զz�������l�����},�RU*�5���Ӑ�cYՉ8=j>�Db��k�s�"s��w���`lc�b-D*�sr��ӅJ�>�����@��Bȫ��~�p�k���[D�b����;�J5��x�q*�vx���}����TP�j����:�/�Zys�w�AH��W���\\J�ĳ�٧�xJ�yE�A^��?��ӗ�5�g��w�١G����^�V�;{ǔ*O#;�\����ߢ;^u��l��a`J���9�7m�@(�7�=I-�Ӈ�<تP� t���{	`1� ϭ51�8U��xˤ(v�_q�8Mw���{�⛭Tvg��G%yL�hOc��j~y��J`i��éqZ)W�89d�tj���ϟ�/*l���.
\��y�eMAA���_�=�ҽ,�v"��ζH $@A��/J�҅���n_�$��"gf�%$q����Mu��f \���=7|1ܭ_�,��:'0��r�qS*�Z�XTd5"���QFL7g���}1��S���h<��$�p���<2{�<l�~��st�Z��h�_~��)�3xK�8�N��@q�?��Xt60T�^�U���c������W�mæW���9�s��䌮פɼ��L�$�eĻ6s(*��A23�M"�~�A(�����7�l"����-�:\��s;��54�p7f���˗�Q޶4��5��"���d)zQ �������0������]��G�?a�b����s�b7\??,����oS��5Ԅ�Zw��4*��|�"O�q���;8�5(�/��ٷ�*++k6���[�,L�k�,�uzQQ$�j��;ojCRFr���ۃ�}�;.�����5~<,(�t��9�۷Ix�+ܣo�/7�8_�@QƈX���҇v��[�5���(�N�]V)�HjN�|� ���KO��z��Ï��W�L~>,|�+�R$�ϯ�53f��ſ��=*����	^�������|�y�G���V:w�^`knnI�������=Ǎ�J� iX����.�\�W��5��X���sc:���J7��ӝ��Ԧ�&w��tb�bW���J�*H �3��N��i{��G�x���ub��Tj���={ ����M��f<\�?���I��mV�I�%o5����?4��O��$E�9��_=�_x>��>����çrD,��꺆����օ�Q�Xm3���8	m�v}��6� A?�Z��S�)��,�?��	�7�祾�u�`V�E_�u��BDn�z��3�����ӄzB�O\�С6�?��	�n��E��L^ǐ��NKE�zw]�_���&��#^��=���i�{��(��!6�h~�՝����ة[-5C�%r��ĊOu�|�����XL2d4��U`���Z�o5t��̤H�I2�9�R��ؽ��ء�/Ӆ.`��yi��C�)�;L��d�H���� ��g[)ie%Y"����}<BO��[j`����4I� k��qVG��/-�������T�h�pR33�6c�3��#HךQ0#W?@��ӛW�e�V�G��bY�jL�u�`����g[a �����tu�Vʇ�솠z���s�H�@�ԭ�p}�e@o՛�z���~|z՟�; �>��Y�2���I�"�?�Wj�]ӗ+]e��]�7�s`��i�OId��8�HF��I�FƥF���+o�W���ϝw�[�����]5�~��ُ�?�"����w��W�W��X�A#=�ǝB��4�TxH�ܜ��t�l��GIz|kvu%g�Ą�! �Lg�����:�#����I������֮�oZz~ŷ�B�������b���&�W�1Q#�R��S�ZɊ�~��J�w���{��P�x_�� �y.击�V�_K��o��J�9s��?�j������ȓ�zָ,G9���@�̘�>v��[�	S�F�, �wGg��G�D�ݏW�T����2�Џ%����G��;��mf���Q?c��p���Z�n�#���F+!�L<ÏH2I7�d�㚠r؝'�I�<M3&�Г�_�&��X�o+2�ǘy�Q�V�ͷo�WdF,�Vh��v��Mft�'����,v'���2�o]���{�:��Fg��m�5u^�7���rq�wg���#E���=Qf�]��f#y9�g�����.�+g���A�����b�a��gyX7*p:�<�t��:`e ��F�} %̺?3lo��u{�z�C�,G��k�G%����R��_n�F ;�a��F^$��Ü��,'{s4!7Ĝ�v��R�?#}��������������TX%��κ�EgOB5FY�~H!ru��_����+`���N',�@V�m]630&l9��їo �$`��Y[�^ͳ��A���������&$��������v3��_k#�\�_$����En��ϫ���1�>�Gx�Z��<���j<��\���O���;������P��0
�.`{��NT����4Q���m�����Uz�/�#�D��n5����3Y=�R5|,4Vm�`K�+���N!�b��.����gӀl�᜜�V�FmJ�Gqeۯ7�	n�}*�_�ig�?'���b�߷�rOIM���6����L�x����٫s�y�'��]�bOL��@W��3q����)�"g�w�3a��ݭU�ݾ���tϻ�b |�iT���Z�/��e,��Ȋ���R�~G��\����&q��3eO|�v���Pi�Z���gB�h��tN���0أo��뫟�>��)8���.��p�jQW�8m���Q�S������o�;ˠ'����NK�?d����O-sMdV�sĲ���GQ_���B`WVjHvL��sӾ��{U[�1�%N#���~�����Xx��[�H߄h��o�M��2O'U]��x}/�~�>#^�P�XH=��P���<�T�][0��l;�:�������VtNu����s�̼�^aѰ�y.b�mT:]O�Z��T�ܵ���t��(.���F���Nh�A%��Ȓ>�}� WJ�郔�p%>q�U	�2=U2LRL�!�$4���`e Ng{J�O1�,�Q,2cR�ӳ�w+���ikaҌ��<bs��k�e����H���V}�{�3�u�.$�0��2�f&p�.\y�$,��cE��T��Z-\������,��~�"�Y�x��tR�j��p�t��e^xu������Ւ`��R���3�n��g	B:����tMx����#��l῰����,�����D��<MN��ݲ����N>4`ē��@��,m�b��p�\��'���E���Rϱ-�p �2�3���r5�qE@�@@�Ê��!�~��lq��<Ȣ���b|�̓W{�P7�d�&��j��u��5١�I��e����Cx����!�g]���p�%��0%� ����k�����]Qb����)�_pPx�"�1f[ٸd�@,&�}���e;���O�q����{Q<<u~2�P�X�h��eЩ^=�c�}B�Z.z�R�Cw�5,ߨi�#��PH	���&�|H~�/*�Kޗ�~�����.6z�������--)����{x���l��%	�"�"����:rr�MI���G�,\2��������ZzfHf<ܭ�麳���$p�:筨b�3,R[P_�:5�w�;9�=,&&�����Tg�)�'$Ʃ� Wp��喎_���j� ���ϜE�B�r��@�p>�ES��W�ƌ�4"�m_���G�#$5o�%�L�w�sg����r��;�� �����YL^O���bl������b%�v{����6�J~�k��<���x;�o��%�}�/�q���.�r��'�Q����L�T��bl�����/���)_�9MB�ډ�Ę$;�//�~	�U�.�譞"F|��N4�u�+%�!2�N�m$zh�ǳ���j}W99�.�<�H���<���J���d��>���@ �j�J$�g+�7�:���p	�H��/q:'&	����Nt�;��-���'�ݻ�ݿm�K�"p������ϲr������7�g'��� ��p3ߎ�yQ�k:����%���`�Y�ED�c�=	�zo^��d��H�����O9X9=���2-��k�JE����y���-j1R�E(�ӣ;i����扊	<T�a�@O��susu�E��ƿ#�\�����&{X�5�MJ5x�9�<?��D��\ �_����^�`?��	dE*��� P�z6#���Y]�YX�<��a��x�kt�����O��ng�����G	�$��2G�4c���s�i{�+�J�u�Ï���u��С�X2S�q��W��~.q>!�
�� /0[���tM�x��_���q�oo/�p� �q����\�g}��ۘ������# %��4U��#��uƦ��ѡ֭��҉BP9�}r��߿㪻ro�+%@�s>Hb-��4X������{��9�	@��̋RI��C�?�M;N"�#�Xq�3�]���T�vVa��a������?�Ӫ����O����	���_���ׯrx��k�X񒳏3�ŵ���kO�����(�:��3�1y ��/��	
�(E�eh�ȗ �tzJ-��,5%c�. �^�pHF�TN�����^�`?{�6�RK�e�%z�۲))�4��t�����L�v��r~���$рa�"��(���J��ad����Z����8g���}�/�'�^�?�C��o��x:(J����	��WE���Jf:�����~�~~�L����Wy*���\�z�������H1MCK�;,�þt�@�/5��h��-��_�M�\����z��Q��3_�gM���щ9ñ���\F��uM]��(�h���I��2��TS��s짿ӄ�6�>����kn��w7��$�4ܰ���Q��7jaMrO�>�P3�E�4������:��P�2OE �I�� �01*��pe�$�6�趹�y闑�J1��Q����h���MMM�ӣ=����.a�Ӄ�"؝�*��i4~$��������s_M�u)
h�N�ȍ�z�z8�??�C��pSFj�k�5=�c��Co�T�x!N��Ύ����������֑?bۉ`�t������ڒ0��.3�;�\�E�Ue��@�u���d��!E��tpe�ܦL�-�+�
�ќG�����@S;�('b�8��n
�������3�eq|�D!�0�Bd��=��+�4����2?����ŝ����E/���>��ys��Y�kʽ��K<� �l�tV�}~���@�A|�i�U��SAj���g�e�n'�ۭw��=P���r�Z���1��{�>�� ���ؼ#!_��.z���`x��ˏ������o��|�a�^1��n�k8a����CG�\�3;��nh�ū�ؤ���0�2�;�njU�X����!M�0������!>�8. ��ڎ���$9=N�š����;��4r�4}�'b�����K��zŻu5��U�]xuwT�K	U[Bm떐j���+I�ˤ���\��<o������<t���V� d*���F^�l�}�ai��*CgU�Y�����ާ�xj���60���[0�OZ��m�+uz[�3>R�5����ۆh2��z���[z~q��Qv,�.��kh��,:B�8�t��@��s�J=�p@��o�g�x�y�	=�t��2�<�]IT��T�+hŶ������]hj$�9i�����O[s��y�I����_a�v����&�_�߽��9>���{�j�3&�QY��@�'�}���t�ފחs'_�׮�ǾU��������6�N6G��#V��2��9�d��@�_��
����,��a���UBey�.���\�6\c�$��{'�}?�kE���>��T5����c�v� ����f���Qi�������z��Y�����K��e��ǌ���Tyg ^Aa��&�G#�o��}�����I�Җ���DW�n�v9�wJ�COs��\�*O@���:ͣ&�XJ�?l:=��&l�Q��:6����ut�>�?0�[��ӽ����oö���E���FZ*te�����aK;�~���?Xh�ۤ�7��}�{:0��T��a��C�2!���F)v[�]xo��)���r���0���x���]gq��b2�q�ՍI&��8N�~���pT�����eD�N�ưLa��M�6�X�R��	�Qڬ�R0n�і-�-�o��:Wx��ϱ�Q*�w�-�v���m�5��mD�9,R�i��p��^���W����m[���oE����������f��	�1�r�V��ű�>���Z�U�+fff_^����\J�]�/lS���_�<�D��5M�.4jx���˹O/-¸[ch�D���Sg~U�v�M!��[�`���t�v�����\�r�h��Ks
�*�4�Gz���v��k8�M������R��o][F!�A�/���_ՠ淣S���z���⏨������vN��ZE��ߪ+�8
J�R.�b��p��� ps[����_���A\24C�'�恾����K�y���ZLB����`��ׯ#�%%?�u?�K���O���\���~�
ÙE��RN��ç����n�0�y>sƐ�N17@�]4 `\���R̜�҃���Zfc�u/���vSJZ��o\>N!NۗH��W��|Ʈc�������3M/��m�<� $:���'8쎊��$����ť���~z�!��Ʈ�Ν�e���Nz�̿@��Irh��c#���`M�x�&� {�������J� �=f&��ܶ|}}�R�
�=�(֣�҇�xD� �}���z�jx��xN\rt�d�������zh���ܾ"nJ�u�]��v�B��아��5��]d^+�Y�w����3��������������99������x<�Ko@o�%դ��Ǟ��R�Gs_wI��$X`6g�-�ǿ�D�$����{]�z7-X��L���pJ�{r��[��#�O�W5��S�G�R��8� U��72���	9���f���3/2s�k��PU�!�j�ǯCO�_'�w�2��-g�٘L4<��wsi|����ؒryTe�퀷�1��Ш��Dtp�<W��(��������Z��p�ଙ��׳]=,����]̙70�[/�!^��^��C�,^�٬:;>{v��:!;��5��`�xǋ<F.�1ZSgv0���u����Ն|��L� ����Q���*�>8�^>%ݕ�;Xw.� ��x��Ħ���T�����2�̓�?pm�b�:�w>��vSS����١�6�w'<�첊�#�"M��E%ؓt��9�����깈i�す������q�E&�N���C܍�8#��.G�].�N�Hb;`Q_aNj�[?��yZ��������Iu��a E�W�wK�v�kdL�F�a�t���3�,16��ۭFd��Һ|z.c�d,���"XX׍d�o��ä �{l5y:=�þ��n\r|�թ䟼Z�$�4r���n���H#��%,�.��P��������wJ��;[�͟w�w�,���n(
�$��ʹ}��Y�(�b�Eđ���ȍ�A�{�"i��r�L��s��+�GE	]�/�'ͪu��=�N�oyG��I>f��1���;��ɹmå�gzѨf����G��"��ӽ�Zz�W1ū+e�dKuY��k���'�����Zu� K ��u���ͭv�9�zݼV����KFW�7/�Z�X%�^^����y� Ko9�a���;oi�)��?����8�����H���)�׻�}k���������?8�|��*�m��2 ^0�d&`��=#�W|�!��j\��ğ(�_W�~�p�'̼����y��~f��cG��י��W�"�#�4�NB�*��NZ=>��)##���I��|e��c7Ap*�	G{k�\�i��&�~/q��9��.<׹�ζ�b]z|giq�yG�`2�;�_�t�HbO�_���� ��y��{o1�h%Bb"�C0���&Ȯ5�������}���M���le�����Z�C�^����K:�U���ܫ���Ѫ嬵���n��>�Cܑ�~�uT�^Cm�:��u�%�gLn���n�����F	%v��6�A�qEA�2���Z��������CA��/�4����W�����`g��^��I�Ű���C��e>i��%b���+�rQv(E���@x����~�����>O]�S~i�Z���-���35Z9b�}�a��Gb��SY��g�p��Ӱ-7�oW���s~������gkD�U ��j����_.����CȺ>�L�/�]���u�M	��H`�
��Q��|�Q�^9����:^�Ð'CL �W��e�5�h(��qz���L���sW+Z��u>����F�o�E����ת�3�`;�I:���a��Nm�C_�F��#ݺ0��T�V���eq���j���~��TX���X�P�:��{��"�T�54�DӍZ�"dYa�Ѫ��ǆBC�����׳x�3	Ww����l�@p���PǥMp++���D�QӜ����l�ߙ��ux��4x ��e׺��@��I�<�����=�F�����\���5r�|	����������.w����ǳi���N�93w���?�U�Ꚑ��ZR~D�:�L�����iK��v.o����Hͅ��$�ι��T��3!�7�7����sj��_�յ.�^W�@<� �Z��� ČJoy2���%TO��]�"���]��7x��o�C�؜�\���̔V�X���.��VS�˳��f���F�Sr|��:J���$KyG��3,@/�'������x��o
rgLI�������Ң^[[���������47���R�� '����;Y�`1-���$�t'��k׃��&9j�u��L�w�9 �6�nKá������� ��5�f���x>i{(Lz�]Z�����"��Q�c0�a�������ʨ|�Yk��me mm%5Ti���������!��d@�,���0��j�p�.�����G�:�?BC�*��~Gy�.�Ԩ�;p ǎS���ow|�Mիq�̙�fK��*��v���O���h{�,��.��fr�}�3W�>L��ė�52�vj����0�ϛ�����w2i�~\��3��Z�Dm���p��ȋ�+~zʜ�	ܜ����2k���9sRI-�k�����b>ztl7Vvʵ�
��;�X&@Κ��=Њ�f)�ܲ ���:}䌏�(�-:��G�Y��Xh՗�p����Ue��g'��9�ߨ��f�k�_���B=�[��V!B�duy�4�v
~qBA��N��:IΜ\���ǘ^s�����'��*������ų�>`���2OW�7ⳬ��w�� \���o�3@7��n��U���������!,�_@OU�-��7�t�>*�8z��q\�r�?"�a��JU]��w55#��.dD��x�D�Z�L�#�k���A�M����c��$L[4oW�j�1���H�4���s:c��!V��K��)���g;��{B4�6���cZ�A����n],;�vh-+ur����a�x�!�,3�Z(񁊫,��cz�U٪��^~�o
d1�QE_?��+$rM�adŗߗ�������8��.C��4�^������g|�2(�"��ө~�o%;����z��5���і��FP�T�E��k�Q�C�>��q��E�\f�;ES�KM1�3�����J��f���9oզ=���7������T��Է�xh�,�*!Uh6�"�>��ˮן �b���/�Πdǹ�������!��g���������Z"�:Y^����gei{h�m�����v��kf��f}yM��@����7�i�1���ʮ���wI�rn�~�o�lm�a$e����?
�~4S}��!���D��L�x��������;��pL���Cu
��áT o��IEA��o7��♀5�����޶�
�83,z�=�>�ap:�i�(��$�u��G��"��y�7��L{�`�=�Ok{s��������o�H����2�S'��IiM�-7��2��O��T��e����}8(�h��W2V#���`��
��e �kmR��E��G8�;�當v�p����D-�7����7\j�b��;)�$l������d��O�"O4L��g��X~A6��4��ĺx5�^��������f��, ��/�*�t�#�:̅6t�3���x����O9L&��^�!&�!���wV@yů|�L��,W߾�;;��*�w����cYnkJ��*N!�4!!���>!���e �M�ؿ�$dWhzֶ�� �~Vb\����n ���(�|j+\~=����&��O�ȷ%��&J0
��/d��7Z�R�r\�&� �IW���W_��r�J%+�%$��d��p�M�����h��� F|���Gџ!a�{�[��8B��{TE=�A� ^@J��H$efe�\��J,O��TspZ�>��\c�Sdn6/^/�F����4�o{$V�Ԧ�2gkV�>�.*�= �`l#�*C�ن�ͣ�~�	��]!�L돐�������3��y��m�܅��Y�4b��8p�;�p��^�hn������s�N����пˢ>}�};����}uA,---8���T�4��?�_����� ��� [�5\���5t�Wq����2��G��?����8�s�SMp�Ђ��Wq�?�B�|[|Ipp�o_�7k���L�V"];��I8h�H��(!�d��������x�BI���YK$+������F���ИڑJHH���jc	b1�Zb��Yq�Z�)�h:���G��}��Ov;�������LRPﭫ}z#��!.�ӳh���*��T��!�[Y�馜T}4;m���vsnhF�r�" E��d�IE��7�K�^��%�=��8e𹳡

���%�r���=�OMM�KH�`}���3���QsSP��i/�:��n�ՙ��#�EL������ �����\L��E����w��_b[�6���Ю�[,�x+Е����c937g�p��n�`2���qrԠ�K�Б~W�����������w�Q�	���ɂ���|	3���D ��z��3�J�^������]9�F�f��l�M�����X�_�ƽrb�N�J5.�P�9@u&��eGG�4UA.ۇ���tl��_A:_m}|���  �F���{ZZ7^�I�BG�.��o�*��Vu(p����ύ�V@��Y� PĎ?jL�A'��g��ot�Ju�'[��waᖢ�o���+(���I�+^� ?�祅�}��7��I��= ��y�t\�ߎw^��">�U"�x5!����j'�5�*A��T�͏&��_�J�������S|�<�3���f�X*2�C|��$%�ff����mU���ܠ���N9qqqvNί��E8�ܡ���
���l��&~!a~O3�7N��+rGCp(�e+��{��2?vZ����+�Y0�����V[m\��<08(t�������֚�4�ͅ���R����W&�|�U�a˷�h��E�~�Rtż��D�L�h�7�Rq�Q߼^�W!������e&��9 �+�-�U���/�L_S_���[ �NM�x�u���7]y��#�/����"��%�=&!�����7�:;��d�㣔FxUd����8q"��oN��z���+w �d)8���'~|~!�U>==���Y�a�RIv�@���[��'~����Y��أ�s��_���#�U!D�0|�c3��W9	�w-M%e���%��Wo����gRy�ܱ�UQV6���r���������(lM����j�e@Br!�S�c��pڵV���SB���8��W��U�O>!���C�X�C���ɺ�������X�-�2i2�|L˚���,nF�r�@�}lc��ae�*1�t�ⴖV�[k�w!�����4=�=���D��|�F��t�cDE2P��k����|㯞�ť=���2=s��7xG�,T�.d�` ��RC#!T/U��C?=��������ݸ�;]�B|6.�ua��G�1%�!��.��<��"3�^1țW��Jݠ��=ɖ��!��B�?g�������e (Va���o[��E遀X�7T�ɬo����{௣��`)'� �,x�:y���ʅ�iK}p��nR�,�~L�ǯiQ���xR��8����g��	{��������OM)���@�~b��=���,|������Mj5�@`J`���|-ZYY���������'M���m��^C��ϟ?},f:� �x@�A��юy�����3����=�K�.����Q���c��;U�Óc�{�GY�T���7�e��� �����f�^M���\y������Z�_Y��p�t�����Z��y��э�"oI���l����pN�p�_|���X�YGA�$8<ܥ��y����X�?|�`��vv�I��k恐�-�˗��[��_`Z���[�e����&�Gȣ,w�R����[]�]�8|����s��� �/>���,pN��ΰ5��"�����O~����W���ȕ�n������|B.8�.t�^2��}u�SVH����I><�!���qf���|��Y��B�qK|�k�cOoo�3��\��������=���A�����=�_be��	�T�\�K�.D js�ܹ�������g�ʟz$���=�q�6Y�yB?���f���r)�J�IV
L��	�����;	_wl(�γF���<3�<�٬>����S�&�4WX�:O˸)iM	��{��R�-�m�o}U�k~R��Ç�	��v:G��6��1Ǝ���$���d�7b�W����fɖ�l���-ڲ#��Å*c팷m��aL�J7�;&��%�%���o
��Y%�4Mݲ��54�����4,֫n*b��'������
:FV�Łu�T��u���>���7�����FNT�4]2�F63ɀ�.��_|B�
=v���3�]\ܧ�3�<��=oL����q��jeR�^a�Ƕ�$�g��˳h�(c��ݛ[�y.R�7�_*d(����1x��\���bLE��bi���y��[�sIڋo����)U�{\��<�D�f�E�����%V�0&q��e���1_�l�s]܄+����F�U|���8m��0�5["��C��Y�=ƷٔvcG1 9���m�X?�U	b�4WB��޻B�E��'ZO^��@֕t9N��7�@�)X&�X���%c&��k��lS�BG�n
�{'�!�����g����ʘ(�v����﬷���h���,�LUl
�jW����>�3�т�0ۮbӧ�C]�%����^������"����G�1�$j��m�%F���k�J�g�޼�y��OW����EW�F^u��A����nҥ��'�q�/,�H	��e�Sh����A���b\�w� ��=	�D)`���$��
�*n�v�}�����0�R���.���^]\��X�`���B��j��$�[wC(�rE0�f�I"���[M)��ö��f�u�M�詒�n�Y���������$�������Q�qb�/~�9X��iwн��Xe�d%$����?5���d�лŹ��i�2�����a+*�0�Ɉ}��������m�0N!Cc��Mх6������6
J�R�������'N|�D�I*__O���m��1��R�z�;z�J6?`��b�v�*M��EMlQ�l�Lٍ���8v���صIٙ[�X?c����@�p��Q�oD�����,�(��-#�;�'	�4��|�g�Ž����8n�/>�~W���o�h��p�j�ߔŪ|WC(%�HBg��Ԍ��tY�v����5�4ֈ�13oI��d$�`5����𲴻�������/-w_C|�s��"#O�9����9ޜ2�9�q���]��u ;躳�ŝ���Nt�- l���#~�V�ze�Z�40�`�>�ⴚZH���p�m���l�)����i4�#|�k����p�!��o��g��1a��D �9hy�eңS�.nv��wo�U��[�*��{����˷��W�$��a}�K�{��D�4DM�}���e��hl�oxb�iN#�9۷�q�J���+�ן�&�
x�q���l�<W�*݃$�~���}����hP��`>P�3��G	��B����L�Q�!�𺬗�_X�t�6�(�����~�;ɒn#,����o��8��K3;�������Klo8�?�������g*[�{zz��[���!J��,Y�oWO(b�a��TPEM��<�
�\[f�)ߎ��̀�����eZubE���/~H������#�z���0��5D�����x�@,�����U�w.��F�Kg�[�V����{�W��.T�]ρ�M�c33���Lμ�0[F�Դ�?��������i�VY=
A�Kr��}��ΰ�ta/F�~S��!=�:��bz�8+⤹c���d��C����p�3�M\o]��6��K�U�l-~�$P&Bˣ��/��Sɰ4d�nڢ��X�"�av�ɥ�DDZ}������o��p�_#�"���z��J�f����Rȋ�g�/�6��*i�T�/Z������?N�;�JL@J�c[��՗�;=��׎�@�v+����X���=nM�	��[/��\eRi�����s��ɐv��R���'�?k������X	�(�����='�z�[�@h8��e�ޫ�k������{��H J�Z���`�$�g����vR��Y�I�{�R&�\~�F[ 'Ġ��_�ب"ek�f��Q����Ge>����3�kp7�ƣ�����-�5�
5�2��}�\.��sED����|���?fg��F�Zi�+;�.JVD����6jn�<(!!Q�_Z�CPr�)�._���y��/,HE|��%E��8S����nU�8��yٛ��;GJ%b�R�4�c.�9���҇W?~̪���Ћ�jl]�p4�G��Zɛl�I�,@�5�`�Evn|��`QG�Cy�Sd��l)�&;�h�����c�<j��`ܧИB�����."R�>��i�o}�}`�h%it�q�e5ʤ)U�is�m�\]P����?�'๫b��5u&�����qǹȜn��o���B�SA���~��hp���V�]0�h2�~�I����g|s�sgQ�@C��P�s�݄�MFXtǝ|7�mm������:P4*�=�}I�2�~��+��$�v}�};��1"��Z������߿������n�������lu���P�ᐳ�{��=�����͝�%-d)�i�T���@b'W���BġutR���D�p H�Ӏ����S���!��[���R<|N�o���y���_�h��:�j�,��A}H�F�4X�����S�N&���k�eG���θ�O��� �-�g*n�����W��%�1l���c及G��ܞ`bٺ��Qz������<v�vke�4	���Fe_�ag�g��e`�q�>4�K{($}�J7����p&����۴�Ý�:�NՋ��M��0�ݧɡ�`z`����Yg{���-��޵�~�.��Y?��ez�7�<�+ڡ�(���T�iݙb��&'�E©���b�U|���������qN���wK���9O��U/H0lv��uᩇu��(�a�>���mnZ��)�
��iQ�'U�`�Ⱦ�%6 �Ң��"L�_&J�KN|���0�)�@�nv���76�g�~���������T��귄3K���v3m ����'t���C�$*����3����jt��x��E��/j�喐H�;����;fs+��.ƈH��O�.p|��d)X��&��1l0�-��􏉔�˟���a?�h�ne6X}d̟{@��8�O���dG�''��%	�(b���M���?�w�vQW�.r����B߭�o�_愗�m�~/t���O�r��
Q �	�x�0�l�~���E�}
B�(�ݷB=ل���a���>!
�C!���u�zD3ږ7,�#�Ӱ�ձ�`�4���Ϧ��������[���ĸ�B��R h��=FZ�����8͍����������uǚ!*FF,*��+ZN����\_��G=ǿx�&��a����6�sq)�D��8V��Ȑe�0?����=�y&����-j�o����>q^����̀�Y���h���}��9������#�ϋ�&=$�*����Qv��3�zw�� ~��>c|�O�ˀ�d�:79+������k���ޫ,�[�뻣dר��@�s�b�o���ې��A%��ג�V>`�0t���eo��:Մ���v_��R �R$�F�_�;2��Gv�`jN�Wz�o�yVu��>��@K����#��n�Ƙ4���/�ijj�����|�ݛc�l��|hI�pL_�+��*0e�RDYKzm��&�us�����-���.�WK+Us?$�dt�T  �;���~�;��2�}����M�54>�TC?��%nk�择�s[3�&�֝$���5 'W]gz���0�SA�J������8�޻�><$2d _��I������+zb�Xch���Z��\V� ��)hG�t���������p�y�ֺO9\��F�{
����&�[P���#`���lC�Z[�m���O9����0d��κ��>ql�H��ah�6���/Ҩ��Ď��֍-jDY��;�]YP����ǚ�s�h%ݏ��1S�AU��d	[�Z��7)�t�	J�vO��4t���$�����������!`���霠� ���B�}`܎�7#@x�#�8������G��7['��l��mؤ���[�"Y����w����ڄ:��}�$�[^;{FHOþגQF+�$���ʎY����ӱ7����5]/}4N���� ��L��d�5pfB�l�߹�3�ZW����PwR���$�W������_������d"C)��#~�\V�|��&3��
~�TvHy٘z�v Z{��Q=���o�	�\��L}N���7�|��87'�Y�����m(f���o��̌��.u9�s��x�	=(%e���Ӓش��XN���a�؊�@F�%,��X�~'|�A$nG�OE���������_���:��=c�j�1�a�8#�S��b�]�
6`��͠-��<_�[d�@�p�I¡@,�y�x��l#��! ���h��W�y�x��q�� ���g&Zc����-(f���K��%�E�(���
���> �_]�5 �j�����6!/Y)��  �˦ԥ�zߠ�-��s���0��s��F�A��]�	����2�9���(<2$�����$�>���#�N9�ܡf�7P|ے^ʬ��t�9DX�o�l�V�a��Y!z;��{d��,��	���<�&�a�,����G�̌�F;�f+�|������W޲��#G��]���£+i��0��mk.������؏�
�w,�Qc2�%Nb�TY�u��xvq�"�-���O`�;N9�$Z2�M��� �PT�x�plZd��U�A��^��@�e��Sy�>�\|4��Z���]������Z��p��¼�%H�k��#�K�#���2���A�;kc���8q"V��Y�Ȥ+ �T@N(`���D�KK��K�
a�<Z�)𒁙z �>ȅ�l�A��
ԋW�O�:?�Q�;k���"X8��7�T��{o�WJ�t�Z\�;Λ��M��ZK3f�ִ���3��if�G�/^��Bzl�U��ev-� ?����p2B!�i�4)큍��_�&!CX�z���o��Gggg�k6?2_~x�lE�#a讫�����Jڥ!����x�Z�(Z��9��g�ːF\�^�N_��߽�ʯ��C4�X�z��F03��\�������*������h/��I�)}S~�uT\��O��D��J��>����Ȑ�n�\�9�X\Z"]��Y�휀	 �A�%���܂���1�+s����
(�E*CP�#*��8b|$���)�`g��<��mpʀy�(�-4׵k��+��k��.L���R1�,�;��ΌV8�4 �ꌋ�n�� ���I=��~c�'�Pw�Cg5��u�6���"�<;1��_ �u����+�ƈϹ�{`���\�!����}%�\|v�ZON� ��4�����%�R���
v��Í��}^^^`EJ,�
E]�x4_���P���
+/u�<�5x���'n�P��A�s�5�X<6�N��Xj���ܥ �t��I���Z��2��}�9>�߱9��B���ZfA�0���M Yg�����㻙C�AM�O����0ֻ!3Q��Y����N���*S�����S�崲Ut�.���xY�]d�h��53�:!>�T�a�ܞe3����0�%�Y���k����m��k��c��ʁ��в-�"��-q�4oP�<{Y��$B-IL�i�o����n��B#�Q{��w�w��6Q̨���:Cat�J��f%W��
}��Cx3=|����V��|(��t�:}\ՙ�0���o�_�fHI�}�n�y�����~�*�:������V��雗���sr;%ԠU�'Ӵ�ݿ�H���g\{lrz�<��rD�W��ݮ�=[sL�l(�?� �.0>>��ɡZ�|=��!��1
`�֗��)J���h���}�	���L�6�jeic���A)w�Β�4�¦���p1x��ՙ��R&|�%,�c-;�����M%���6���#l��t6u�lC���ek��ѨZF������:tsI���
��g!�s��`���3/䗆
�r�wtw�H��`~�(蚾𜘜�E���dw�JI��Ɇ ���`��S�K��21$��"�+�+s�l�L�1�"���7ϐw��<3�|�PS��I��38�����δ�6�w�E������]IV\x�`�dmQ!�1�n���X�N������x��x���ϊ&�CI��Pz~�A�ON�͇	RE8�&���Z�o菞�څ�ʩ���ve�/n�OAW�WԘ���j|wo�ﴥSN���MK>�>���ou���G�WdN^��`a�N�Ğ�b�D�l\��b䃨���]���Q$����˻eu����콒��b��U���4�$�I�bUt��?p���_��,V���Ջ��6��1���.jhb�¹�������g�+��Q|z�D#8�G�n��}F�����_�\� �HI
�x%���'s�~��a%�
�FW�N�U� .(v� �$�yxZQ�=ub�£}�q���%���b���d��E6ZZ�ܘb��keӛ�ng��,,(wt54hzdJ�7&���E��w`�8u�C� �h���מ�� �����uz�l��c8�@˓G�8���Ӕ��8�"��oq�<�9-�v��$J&���F��k�U��|��������v$�vE�HR�,�![~��R�;:\�zj��v�a��ާ�
GA���	8B��W�ѣ�V��L��8w��y!���8��%\A͎r3�>f���{|^4�L�" ���w��/`	����|��U?��Fœ(X�l�F�/�q��z�q������'����K��v�!U�/���Lv��)�^#����_��X��� O:�F���uT��@|�� @����S�D[�h��Zo�Ǳ�J5��6~а��Q���= �`]�N�����.���y�䊸���u�kO�'w*��g�ߦL��O24Ԯ"��ԣȁM�Y� (`�_����h�!3��c��=���'�D.�zSa�b�7���Y�l�2.�_9I� ��I��g��(wo_�o+z��2hR��ө�U$f��@��Ǫ�\ǜ�^�V��}��f��]oAu�O���$�73@ɰi������4c�5�D0�`֛�>�8���`WUU�e=�] ~t?s|J�\�q?���D�������f9��1#C������|�����	Hq����i����U*�����Qsx �[���':m�Y�����D��1�,ug�q�K�����6��F��Z��y�/����n'� ww�b�l��6����[ �QFO.�#�M��w*�	�q#S���F(�v,���X~�U��6cĆ[y�v����9k�q�h�ڱ	�)_�2^{Ӝ��vŨ���Sm�̌Y�9 �Tj������؆际ezI���_�����A@1錘~��/��Y�2Fg��וme���|1Ԗtܹ8�+���~p���Ҧ";_x�T���Ė��R������*�W�&���PCOI]�.iH=����п� �V�Vi ����o�-ӹ�X~:����J�(@|	"� F�j��D�Yn��AD.@�}6��;��Sv$��0�@�IݧM}��f�~���ie�ˉ��v�ӯ6S	*B����6��3bQ>>;��/Yo��טlQuwO4־��-�-O��݂���<����~Qfwɩ�lB ]6�W��%�}��<$�4V�_o��o�{��i婹�V��D�:_�Qu�Tݤ:j B�+EΦ�����W��LA.>�$����v��8�r���0���ߵ8D��@R�}r���g.�~~��#����tu��7'�E��ͲHIq
����>.+�Pa�Qq���ގb��b�8�cd�co� A�#lc���ґ��Ȯ��r�T�1��{O�ಢgZ��*2d�F���ֹD����4��a(�,ҋb�K�5��R�v��=�w���|v�&�e��aG�O�1���s`�����������	���d6�W��4���:f\4SWY�.��E�5]n�]Pߵv,%� ʨ[c�kWQ%�9 ����l4�rbf��1�bڼ�A,[�FuTτ�.��,ԙ^����� .>��lg�dB^G�V";#G=�J��	 ���aLZ�Z#f��W���T�o2�����0���TN���n
ylY~t���0��4��'�[f����֥cOE��(���OCCn��,sM�R�y���	�V����h���0�	�T����Ûw||j'�Ͷe�D ���O��O������N}�oRR�$��~�;�1�>�>���r�~�����L�WW>�y8l»G���%%�J���!&��+8~����	�+W�(qϾ6+S#r<vWW0/np5�n� e��_�b[&�	��#��=c��N��'w!�4f������`�H�@��kh%H��Ga��}9t.彻сT�V�˷���n����t�9�cv/�S��i�	z- /�F"�9��j�R�]�T�_ff�B���?	�£m,Oa.))�GO9�-p��_kQ�Q���}ؓ�AI��f[p��%�7�K�P�z֥ގ����b��8B����=���'�~p�y�B�}f ��e�S�-ش%e���.�|���cM]�æq�KZ(����\���}7�Ě��2�� z����S �]�GFV*��h t>�=��e�gI�<�k��?#�oΡc����}�6�F4�w�L"� �'�5�(N���Z��Y���Ŝ��� ���<R�<�M����yh��ո>�,�����ct�:��w�����ߞ�����e��q��SQ����k�Ӽ#u4Y/�����C��!�&w��˜�wV~H>n݈sk'Dt�n�a��3���1Ş���;5�%��q�ysl[Nc+V�T
�j@GO��"�	p����$���x����q��8��Jp�,K48��}��]��c�c���(�T;�Zذ�cHܥ�f�ۈ���	;�Ɉ�6�v��g~d����]0ŏ��TP�+�i��<�J���`���9UTT)n����ނx��l��tދ�BZ��^�_wˍ�Ƙ�i\�5���X�j��q�/���4�������և�����e�%%wq�b�*c ���x���=Gm�Ej��я�˺�lj����T9�k�R�"��~��A/���K�¶eV&^%���L�vbQt��l�d���KD�kՇ�fF��w�a�����TA�T蚵=�|_Z����y�{� &���/?l�օ5����F����x	BB�cIp���1�A��Qm��ؿv����y����5�NQ}�W�7�؄o���O��qp���j�<���4�hJV�����_�?�:�/�@�;�m;��x��gTN�6b����HJ�L5�y��$��bk��������=淎��K���z�ؿ���~S��rׂz��/�Mk��Y���_]��nZke��@�Uo�?�V����ҵ���8cV�l:O8}ʉ36l) �tY�Wf�^��Ԫ��Ӭ�FP��x�ۍd�|ч��t�/Ӧ�0�ٷɰ�ҁ�ݲ�/��j���?���|��R�h��;����7��m����'�'���a��|Xp�;��2�^�D�br����W��'0_�L�Ԭ-4�߳ƏE�n��r�:��xO)l�Ma�6TsHw�ڢ�ق�Pt�j��p�5D�/�k��ˣ��)j��_M�c;D�&�G?��,�Wۨ�H̞#�r7���$�r�Et%˛w"G޾|�RUm+  �(�ƀH��X����e�#�i�/���aa�0I�$��,ǋ�sJrӦ$!�y���g�N?$m���U�lE���꫊�;�s�J����d%��䍶��Y�w.��Ά�l��m��#�M�t�<h$i?-^���G�JSl��/\K;�!aZ-��aG7�;0¾��2oN~���z^ �GJ��ޗ�<7�vj�Ν��
�9�Mڋ��M�F,��&�����4z�E���*��������]%H��|��Q}D�I�[���Cn-Ն&�4ern-���v�Cu>*��3��g�.m��:34{/+o��yv�k����xh#pp��8p`�ZGO�W'{v<ʰ�?�����v�pIR�r�d���ˎ��U���y���9��dCN��LB:EI�z/]H0^����V�,��O���n�F���x��G!%`(��:6���aL��L��K��`��s@k����zo���щ���ׅ5��	�9}d)/�fG^�{'�39+�+x<Y}bp�mU55��.Vf}��Pf=E�0�G"���N�>��x����:;G�^q���Ge[���fB��m�K�ZG>d��w��?yd���L��/y4��ϟ*�:�>!�SOYީy�K��	����� 6I�z�Kxm��נO�90䥔u�|�/�]�AH��(?ݧ���U~_K�P��+Z��mK7�L'ߞs٨g��C*�'�+	�n�<��#�>hPx�l�|І�W�_"��ذ^��4�����un��O��宾����x�˗ٮŹS�ʩ��Q&ݩ�n�g�3����~���A-���Pߛ!qe��j�
b�ظ��!�n����7��w���`hY�@�g_]M�2b)Fv��}뙕]���:^���O���p�$�5� �F�����j�Nr<ʼ�36{�lGa{"��I�U��]��֋�՞9�~C���\��a����M�t-|��	�ƾ\m~�~UQ�?+���a�ѹ��I�>s<��NA�V1&�Y�hhe]���!��ϟ�dv&Y��%�]�E,�	��h��V��%p#������ l�2Q֞N�vfo�`��{x��᪤�<{[l������wd����ܘ
 ��#Z�"��	O2� G�>�o��,��n�v~�+���$&p���f�c���e�+\Vo,C��)r���X�ip�mo�/�wl�����ϑ��:�Ρe�`vp�J�Fo�a�û1�KjV�jv6�ua0�4}f"��Y�(~h74��8�{�	��YJ4��ҫܻ���*f�`���Sl+dQ� ��?�Vv�m_��D������G��S�cL5_�Q	��;h��2�j��yjBl�o� "I�@�T���׌�;u� )�VK�n�Ȉ�k5��+�C
�
a|f�ټ��M`p�ofR��Q�f�vr���X���A����_�A� qn@�������8��fb�x�;lXB�S�'�>&G�����I1�,[���_�!����(6�,��N���B]��ů7�g�c�j���vr�+������? p�9���GL{Wp�?���y�.SG�~tgn(��q-2n~K��-��B�ª4!a��>���� %��\]��u�]��b���5�M	p�4���뫀����j'�V��j���p����\�Oλ�w���$GL�Sy �B��K�{��>�2��s�h�:4��T����3��hEm4�����~�9�%^�y����b�.����*5�w��]��]���z-
 ��U~�I�z��.�r`A"q]jM=1���}��,�[��M�gY*��zQ����ռ����::Z�����Ʈ**'6�73q�1)�a"�ۈ�fT_@@��@I��ޭ^C�&F�gX Y��NыV��v�5)�i.�j=!���O�z���/�����4�j�3Cc}}閘���ϣ��k����؂�ǟBA����ď�L�?͎��1i�:��|p-��t��=�~)H��U�W��K=�'�t���%���y�R�������d��O}�E_�gr�F|>�����q�PMe��p�" h�i�ET@J@zD�(M�"�)R�Q%4
R�H��:��@�&�B��E�����׷V�JH�9g���]Ͼ��熓��G�;9kn�u��%U��V+M(mo�t��-�V^S)�;	�}����o*Av!�
��� ��!`��M������G5��N�a����C���=��ֵq@jn��DII7��Ve]ō̚{�8��r����J�l¨{ug����#���<2>�>�����x�1"��|J�5���`B?�=�>���3���^�U%ە��dz�G1��~�YOKnU tU��-��׬ͯO��?ؘ��z��e�{���TZ���'/�V;�f�]}{i�������\���:���/_��+Z���a�l�9߽�p9���܍�9փۏlՔ^*8�����7C����&���*=���c��B��\�����5��ɘ`W��翸yms��&o�?A�z����Ip�MݛZ0��(�+��f�Jk���u���[���n������'9��M�<�.����\;ē�(tF[��6��ԴE*)��%*�m��kY���y����{�:V�6�V�å��i�4�.Ch�W!Č�3�I:�Mn^�ǻ8J*_��*�)��o��g�=�����T�Bki!6��׼�0b� x��;$�zf�Փ*�7S4�_�IoxZ�o2`�*;p\GCb�t��h�}�j�5�b��̋���o�������g�6��/�(dm���m�]*��_.^yC�]�.�<Q��^?�2�-`� ��$�u��W������n�����g���ߗ΁�a>s�"��Q�!6PDPg`�^�
9G�yM1�"�!7O��P�1T��H��J0�Z?�"m$��z�3�bR�n���Z�?i\�vi��u���KNp;�N���8>��!{�`C�� m+���p���Ђ�U���d��p�#_�,D�r�Ƨ�oe���D/(9;�1om��0V/��3��/�����p�ݧ�f��3<��C���� syb�xT�e��d�
�
yf�E�_y|�Nb��CF�K1T[G^�ϛ����!�&kg��5�G����P����Pjv�L,�����<)�>�`(�h����C���+��x��8b�؋��D`�R�:#�z��1-�YaY�[��D��*�!*��J�S�	I�����!�m9� ���Ye���������_+Z0)�[蘃��V��L&�I�Q'�,|)�X#V��&%�r+��-�{��Өop�5ߏ)~HK��]��\�ih���?vg,ֆ�!o�����g����{�쐗wԭ�΄/���OM���#wj�G����bȾe�3L5M@V�IF�}:$@=r�N(O��
W�I]r!�,w)8����|���v")Ο8gk��S狙$�K�3�3�l�@�LOjZ�����%�^�h�&f���� �q���Ew��X�?�� �^�l~������~����G[q3ŷ�;����T�l�|r�y�}p� �
�`�f��zZ 2�M�m0S�籩�}T����DP�7�{������tZ�\��+�Km6�!TjM�`�s���Q�a:�$�jz��K�h|Iϙ�+���$z��$c�?�[�k�����ݻ3q�qk�ݡ�B����]@?~����p���������^m����d}Q��;[�;��1u8M̢�k���.�ढ़��LO>ë���?Q>K��BFl�\�RJcq�x� 1j�K{5��~*\��FT����ˉR�����75��2^�#I۵����*y�u�ȫ�s���Kc�Z�6����~ ��y�AT(�:�U�-(܂�n�#�� ���zw6Y�at�0��Ҋ�������Ƀ�JW7�	���6�r��k�y��>;�(c���֒R;�gv"���f;zB��r"��3�~���k�>�Ec��=Qx��*+@;�eφb��Mx?�q�U�t��ĕ��vqV�'JK�-N� ���H�����ّ���	[-��?Wݐ�s�H��h�9��B�8���FN"���<��W�)6���e�����]Ρ'��VG"]r-��zfanZ���3'��R���9e�A�p�K�F�x/`�eJ|Y{u���^��r��KiGs����l'��e4y��q�Æ�f��Z�V/zG\()QN�?��x@���k	���?{�d�6�`z���B8�G�ȡ� �$ٴ�1r!�]=P�s��LX��P���)�6�£m�?�6�+��2�֬޹C
�N���QpI~�Qi�'*�\ښ��)�02��YO���3�`�{���(g�o�N*ެ�$�K�Eh#$A+A�����4�%��ŋ������N��;���b	O���3NQ�^V%�U)זҠ��O�#hMg��5���T�u���N�ѱ��E>8����Y��|f4*��}����P{�ߥ�$���<��<3;{'��x��eDΩ73��ͯ[����sU.�G^n���}9qXڑL2���7���)]�|��+z�4p�Tsm���Lh�Uѵ��yy��� ��!T�nU�ey�౷=�M?���LĂv�B9/��h��nلo��T{SQ�?�n��eo\����cA�l���5�O{�F��(X�_	��y�%\�r��|�qT��w��T�1�i+v�xX>c�rf'S(z��ό���:\�l�M"N�l!�+�n�q]�%g��~��o\A��ǩX� 4��Ў�R���.w �^� �ٍf84��F#���,!W��t-�&��t^����*��mHL�C�w����$3C��r��yG�x-B������#�Ew��U:�T��gpi^@	�+?h��}�b"�t)WZ�N-�>��"�Ɂj���VaҎ����~�k���r��������G�o$;�8�r��*��tҳ�l\T.�t�q�_�q��bHc�<��K��d��4*�Tׇ������@5���r�,vk�Bb�@�W�[�G�Z�C��O��6z��� �	X�xP�{�!�?}&'���8g���8���`�j�c�LR=h�[���ʨ�j�B1jv�x�[�[G;4F%�Qʪ`:3��D|�b��XRTM���q�����J��/�#B�� ��>�K�cS-,0��z_uv\,}0�H�6�E���D�-��w�ޜ6#�w!�+4��4����6�
u+1���~�)��r��=� ����5ggni 1�|��sJ��f]�`1;�V�>�#� �hx���y������;�[��9�����������]�hk�a"t�R�m��v/3]o4�]�ʹ(�!��V��3�=�������*q���}���礐��r'f"6G����K{(��N�gA�2z��e4M{9>+��nk#��dP�R��x7P^��g��X_w�@>\[-��4��.
Fs]����Y�i
7%Ӌ��h��>����"��uo{'�����a�+���A��e�jX�Y_pr{��l�%�t@*�4}�̪a�t��K�~��EǲS���<���iw��x���+&#���
4�[^�8��B�.չ軝��=5�ǭ��BW�^8D?n�wSݶ�������VW�bՅha���]���x���cP�µR�B原mE6��>z3xS�^�%3��:�S�>��:�A�g �mL�ܟA�я�G������6��Ӧ�C��h;�?�����B]ѻτf�Ue��kX��h�F\Eb{�����^Ő�����%��Q����_ԩW�qI���,��v{UY���3�|��R�f\z*�UR
�"�{�I6c7��'�,N�mՐR���Ԑ����A+,ݐi��O�-�}9�P〩�+�;��zu��l��{p��h�@?�7��q[,x��!Z~J�~S����
s��8?��͎�t��ȯwt��v����}We�uL�v��3H|}� �9��3���7���1��r����А�� xɂ!}��]��=!RI�U�E~|35��E�}s^p�LY��в~��f��5���uE��ř����n���Z���v.��v[έ+ږ�/���D�{��ٟ�O6Psl)r.MR�|�}�Q�������-�&2�4�=��M�ϛUڄ��-��!��+_@��`c->wD�^,�KL3����=p[�t�?m9�s �H�ǮeV�J)�.�]�l [m$�J�N���_D��\��j�`2�4��'��.�`���|^�/.����|�b�A�`�'�B��w�ƌq7W�v @���O���ہ�n�QXL?��ϲ�UYYY���p �yw�9��O��Q����^U�� 11�������<����e}F}�cI��un��V�5�X��/�B�C��o9h�ֈ[�p4��++���tdY=��(����i�c"0�iA����>�r!�Oo����^��.#�c��H��E�A(�k_�D�A� �����7*} kaR�)�.�$�{�������/V�꣕��Y��c��ҼDZ�E�B)�a?|Xw���E]]]LN�]���}�)���b��M��ST{x�4;&�T�׎�џ�Kߎ�ݦ��Z)i�]Xӕ%�7ӕ"U�
��Iʝ��$�B���4�j�������US�g-�-�������_X�_h?\�Y�$X�H��;gx*ul@ʔ�6��ٷ�a���0 ��aR	� G���B��-��BfL��6�������^0���u�	�?�a��9?���9����-�!�\�S��!��5��!��O{�X伔У(�4�V!�Kbs�}����Y��)���Wx��ߗOn ���s������%l�>�KBSz#1�BF��9��~��H����e��d��l� �C�-1���hx�a�����]60���|w�q���l~>�F��_�Mn�P�������4'�\���cO��*Mf�C"d@$��3��E� �'L^��-�u��5��d2y�RO��X���o�T�@���5:����-�T��Q�2D94�d`����e��,w�62����vA�A�R^�/�� nE���Sq�i����m��,2j�~��d��\�
�63��u����:"7�������ʭ��䳲�E��Y�6�+�Xr�^�7�O�>״'�y"����tvC�>j�^���/��ᜪ��!�-5�O>��eY ���Sp~��~�{����u���OT���ֶ��X���-|A��Bq�_�3B�k�ٿ^~QT�[@M!|��
zz���2a�eX%0BUZ`LB-?��[YX���ބ�r���EB�8�����k6}���kw�q���v7�f��I* �5 ��L�;p�i#�J>�[��6���J;���_Ó,�#l(5ů̠6~�ş
�
r�&��2�%�S,��E��R
�|9ƘoYy �R+�,7~�5��þQ�}(a��I�1 y���x��hyl?�(jU#��� �\BJn�+^�P�T�*����~�I�L�6�El��G���	��c���:ƃ�Қ1������w�c޿�ɝ��|��mA8�a0�w��� *�+�4�y7�#��^�������w̒~�y����xNC~��7������3���:?C�b �2 �2����7jT��pP�F���\�{ 52 �{��fv*�vt[��	S7�\��D���M^x e,����X���u���4ސ�9�qW�� �Xs�! }�te�+\`g/�{�32.����h�BF��W����+^7w�7��Ҁ��d\����V�$`���m& ��A�b�"�u)g֭��z\��+��.!�y���Es�$�H�K�yu�Ŏy��p"�HⓁy��<�x�$b��/v��.�q�hR�v"��n�t�qT�H�[g�a���6�ZB'0S��Ư���!�xaސ&^�[�('�0;�+)m/��3���`�@�,��1 ����N�ǭ:��^4�	'H���'i��X��k��I�3̔Mj"�/�ȞA��x�ͩOB��G��'7j ��U�(�M��� q�^!`|M���4�Wp��|�Kf�lnmI-�}U�SY/F�9�����A	�$�[��^/�.D�B3�����_��hw�N��8w������nj��v��9�?�M���=��F���L�jC�>�εA��	�-+��S/�ݢ����^^s3�6���v`մ�(4c5�d�%3�?9�4�r���C�ӮC�.e-NKK��$�hXs d�y�ٜPƾW�~˨@�N�h��,�
yZT�}L�w��>��o�R�Y�9����/@��Sh�BlPW(�����L���2�^@����fdW��/�a��½q|>
b��I����I���'�a 0HS�����Ò��vN�gH���=�q�����A�܎k�Q�Mv+%��ꓓ������a�u|v�����g���k�����[EE�O�Sw���EF&V���� �o��")N����|V�����R	�{�A�6��G�����y'�-l`��na[x ��,��	�{��s�
�����&YX��:,q���#T-h�^�s}��̤�P��Ċ+�:+W�޿7(F�\���ΪQ*�awo�ƿԼ�����k˝|��+_L���3�F�8^Rf�(`�p|;�Y�u�J�!)I��plw%��g6���TTkov�(�#��~XmL�NJ�G��t�p��y��Mu5��C��K���N<�Kx�`�|�Y�����m�J�]`��p�+�m�jc	`��e+���S!\�)�F(�@A���f�6+��if�M�;s"�/y����\���g+?�n��������sDF��u��ĲY�?u�
���;"!qVܢ\�2x�����?�Q�3��؍��|��PYT�0�N��l���r��'ۼ�?�@���%d�v��ۈ�:��Ӛ����Mj3�gK�ڗ��-%�8����I47����\��<��7��#b����8��yc������P*:u���x�F~D�}��2�H�˺K���e��
.	��\��AS�d_A����"�A�����ɹ�t��m������"�R��>���7�����!~�@�.DN!������-<���g@|f��?��=��^�A���ց\�j��RA'-�@J�� �%C�q�k���E!z^=�A�{{�zN��S���* \!��)x��sE��k�G
hν�݇���V_���������c��@퀐Dxs:H�c�N>|�eB�нp�e�rrG��$�\�v�^���ѓ�w��5`f4��!"7���?̸�#�������1
K,��6���'�_JژȨ������08(l��aˠ��!��G2 Mŝ=�=O���7�;�f׻��6*׳��W���5������l(f6����up�Q�e,I�q��9��҈h��]��}�4n�A��R��G��BmRY���� �[-�C�#�%W�M{օ���=M����Ƕ������:�dg��\�i�؞\ޮ#��������u��׋�n�3n�_�?5�:�ަ���6�h�����yno�x���jeUU]
���P�A�3��'�<�&m�
�I�hrOnm,3G�T���rMq����� ���3�<�� ��۬��᷵X���9��t���K��~�7�����T��sss�N�&�O�wz���޿�W`��r�E�Ţ#��*��P�%���T#S�<NcK$�'@�e���� �����̥U!��[[	ݔ?�z�pR�d~��+_�(D�͹Xa?�9���B�����#� g�Y�b�#�(��y"�E�e��^gQ�F�E�����߈$\4H=����su	��*�أ=w��py�Vm�k�{�0(�9]MM��^E���5��q6@�s���N�%Ҝd�4!c�;��)����"q�jr8�HH<VX�L���8M,+�u?'�0�;�aP�����qpPq$l���8Vˑ�5�Эi��5��|�AMI�(���2� �& iv 5{��7�t)X���y�_��6��if�>�����Yg C��Վ��R��?�:�
.�Oy��q�(��U��R�S�
�C�l��&��^y�ÿ��D7G듅~1\G�����1�RK����4��1��磼晄�j%BJ�H�+u����=���3�C��0�����������_��p�	��KI/�ݩ�1�ޘ��+_�����V�pTa*�w�6�)��7�y/ou#J��!��mK���F�PA���j�AJ,H���l7wZdS�Y�B�%
��^D @dQqn�p�����jP��e]w�Ӭ~����dr�L<)$��Q�O+t�ԇ>y�����M���&��� �ޝ���7>&��
&�����Pl-�������H���Z�͓m]w])�`��A��T9��)�U� VAk�mf��~@0I; wg�Ơ,��2.A��y��	��4υRh��J��H�V��lӭ���ʷ��'�B��F�d4�wIjE$)H �jh�z����	F^r�^�'�Դ��4vp��F�EE��y�\0��G��y	�X��8z��W��[��P�� �)�`�D,�z!خdx
�7�p��a�
|3���D�; �҇��H-$
�JWX?a���Y�sT�W�e�(�R�ʛ�4׮$q	#�q�����gH��\�~o�qP���y��P�)�K���5�P�p�)1+u?�4Uj�t��\���UaY3�^��q4�W�N�wjkw�=�r�<.h��(l���|��F��;k��b�'~�"S������e.��@z]bS$����G>����.Iqs:�)
-UG8#nS1`��k:�sE7��6�?���W.�
)J�[��4�E��?')�ut���[)����>,����&�i툼���y�+Da��HR��b���+ ��쒹\f6:��1d�6dF����0]�_
K=y�G������l�����>��o���&���B�C�3J��J���\�V ��s\w˪����C���:3Ǒ\CS�Dl�A'���۠�
{��x��0�X:\I�3J�"鴲���r�K񏂆�@���q]=���ӳ�����0j\�+�bN8�"��ʤC�+hc�q����H�D�Ir��;z�?hDm&��7?�"!Y��^%P��}��f/k.q���7^�r�jw1�7�����ZSAvI�ˡ���u_������BQ0�bx��MNb4,�Aԛ�X�%a軃睻��p�9q�n��	�<���1�i����k�9��S;=��	������5U]-�����&��^�� �t����'t�c΍]å��'e���Z�>?�pl�u��t�V�.�G�ܞ��O����|U,V����$s)q��Wj\_���pV���dڬ�^�`�+�n~XH��? �ܾq�ެ�B�`_w��!ו_B�0�t�����
��)���Q��!k�����vK�h���_�R�Jb���>��ʵ�[�u��\݇�l��^��C���4I���n���7iQ�����������0H�J�����l��-0&��<����BM~�$/ e_��U��b:RٔT��Zn�k���5��/]ztTR�}��,=�q��o��m���	��=y�ߓ�ݏc�	+�L^���3oݺ�F��^����3L���A��X�(K��� ?����:YA��i��5�ߌDZ�^@��Y� �+�
���eo�|0���@��n�����u%���_��_���[�3��JX��M�Ł%�7��d4�,���hޑ%��h�����8�e�C(������tN��e��Ug��W`d=h~�?6�ԈJ2��!��a�&���g�k-`e9V�r�5_?��j�}�2�`����4��D�/掏8���%��93��m�@��R'�����6?`��_,+o�q�+W2�K�-��{�Z]�CE�s��d�4ʹ[e5�&bDG ��M�mw��/�>ǀA�Nɨ��	,L���������.H�{�_9p�i�j�ہ�$�(o�x�᧡�3�k����%�
ֻV�ü�w���rT��)(R_�; ��jAl	��g��N�a��������,���Mzep&q*�����ޗ��Ɂ�ot|�����6ߛ���]^�ԙ$ф�������@U^f�0-r%��B�#<xP�=T�*�C`�\���2ʊ�9�1�������mf8�Z���K��i��������	�����{[Mj�hV��3�(fe�����1��7��5o ��bWݗB������e��&_{��������`��<���$�W*KK����#�r����N6??7f��X�IkȐ��;~s��l����,�����O댎��`����P�	i:��x���-���O�=z�i������h����
�
�ɜ'�'�Å���ǻ��d&,���.���Y�q���Y�ה� �H���FC�r���]}%.�K`dO�ԩ��Oi�{��p߱B��=���	����s2��V�`�/���:�g4G��礝(�vHd�y�*�q�Ю
^�v�����)M')��7ov�d
�	�nH��g�l8t �N?$O� ���'�E%.#��s��� �}1 ���z�o�9��C/�"�����Z�k����\N��|�,,26�$l�<Q���;,�!��Q�KƦ����0��h�h2p �AQ_!߽{�o;�O*��zg�ц#`�B���r/��9��z�t�WES�ޢO�����C���c��PkđB��Q����k���"��44�k�7N�����R��Zj���,��H��9�J.^I�\]��e�?�5������{�m��·�$Rx�b�s"�.�x�a�׮q1��5�~+��lR�*7�9�Pp�F�=N#��e�6�~`S���4|,�%����*3k0D�KE�d^��V_YXX�h���dY���RSS�aHW�Bh+K��y����@!E�'6��]iJ8~�6�haO�y�{�eεht~zPܣ��8.�r��_`�yKN/� �ٜ�./��:\j�E�}Y4��k-�[�$Eû� Kw�c��K�X<��T;��)`�fP{����-11���a����n�_.�	����w8N+w/D�;.f��׾t�7�㘟�o�t�7�>�z�oj-���`�˃�,gϞmX�D)�u��x���1�Q4��1�idcχ�1~eE��,1$��_����JC�)_����d	]g�)Tn�(#|��} ~��E�ő2۟Vg)����ô�\�(^_��p�)�Ժ��|X�hSt=¼ġ��|cu��U?vyF�p��]���#bbb�m����7�Ǽ��b"a)��5�m��l��]��u..H��)_����yƖ�v����nMvc��-�Nq[���d�ޣ-;-������L��bb��ZO�iL<����`���c5�7�O�W"��'�.���96?s����hx�[4;���m>� o�����L$�[�?='�4v}��"�,?]�G�9(&�"�]���uW��T�XA9����}�f˧_��\����<���M�x���k��\����d�ג0;���Ib\�*���ݜ�C(�o4�,����[���,�[� �Q���|P�{����z���v�<`ӛ�H^�m�5;���~5ntD�ݝ�:�QY�=�	�
x�\y��@��D+�u��T�@?�ԞX�t��\���>+!�5Hw�*ފ~�$F6������>���Lv��>�������͇�{�H$��]��S*�Jv�m���������2DS���dM�z�{�8���5�){P
�?=x!2�.��1��7T{��+�w��qʐ��7�-w-�N�p�@dS��^�
\7�7d�U���,�ί�	L��m.<Qr�A^�Se�A��k�����8��{,�U�h����#N�g#�Et�S��2����Z�-�;��H
T+xى�Fzn�h�l�&�U��f���ac�y�+#UR폸1Y�U���WU�%^�W��+s�/9�9�/ޘTc2�|�Q���Ψl����?b��Ț%�6v��蒨Qa�̰S$��W�{G�n���l�)��5���5R���v��z6tK	�g>���h�P"0���-�}ٍ���Ak{������A+���>����Q����M��-�_O�Ꮜ�4� _/�z��T��޴���OC�d��{{Tȟ/i�M(�0m]����H#?�[�M�ʕ+�x�Acdn�G�vt��}�5�)2�1;뚧�,�U�*�H��2�(����g�RǊ��!=��;{�Z�`�>��4Bq��V��� �����jx.�0r��ԛ�"!סpӇ�R!��lJ�rW@�� �ݴ
�la�je�0�xtR,ˢv&��+��`��q�F��n�b[7%�[��w�����?t��h)~ut��4�$��_,��+D�K�;�>�Qe�5r���{G�I�-�'�D`���"����/���B����C��~s�4TL�-��o��ۏm�aS�����l�E=:��-��'o
�"���[89�aZ0��u�Ɓ��2�|�a�ϾRȀ���C4&Yٹ�$$������:���(���M7���9��ʯִa>�������O�d
�����rKm�S~{����>�?$t�!B�C��6���+��ՙ��:��WlZ�_�������9j�M:�(H|ޕP`r^yS��/�n�� �n����.s�������n[I3�'B��Қ��ɥ�Ʈ7��(�iT�t��_wp�q]l��!c��L+m�T��%ٰ=��C��_=I�gQ�i11�h�U��0�F	q�����4(:�^QjǄ	�����TJ�(E�k�z�X�A0������S͢!���j��B�����<V�/rdB��gd�������ƺ�ZFdUՊҜ;�1�f���V�95 �(�t����a-p�l� ��A�e� ��@�Rh21�Yi�J1����s�:6-��E%�+
��vIT�:�C'�<>����p�$�#h?\�6�����M[�OT�L�-�1���M�>�Si/Ɏ7�O��	2�W�]�1��uhr�0B�_������S�Z_�Z�/KI�B���J������w��"�͏<���t���@���Fy��6����2
ԫ8�������*U��n�Xz�07��hB�E鏿����B���z^(������ẅ��� ��Pc�5ʣFC
��@\���">�'7+�A�F ��H��[X9fP��wi�6���
E����!��=�{ �?eB����s��Y)nG\.��S������Iy�fUk�)4���7��uq5<N���~����u���Ic�{+N�&V�~�?˄�gQ1�@G�T�WgMM�ݏ[Y��ԫ)�}ς����\�7��`'�4)g�����89���[ڊ�R<h� �7��)?�R ��?���}	�V���2���f�n%VyD|�px|��b�Y�����-�lp�����x���7�5^��j�ߥ�a�A���M�%��um}��F�qS0f����L`n���e���_,֮�eP�����c1���?�tS�O=u�+7kiu��(���J����qv�%W�Oo��1N��408���i�5Q��ӄc)�x��v�[1��=���@�$��I�ݻ�X����S@i�26����������ka��Ffrŵgx�F0�Xf�S��7n�.�?z8�t���f�� �ū�7���/0+�~�	�6!a�-	��}�v�S��ՙ��f����D'\5h�l�h�w�F���]�P�7�Zi��Rd�UpYt"��K�? ����G�Q��)gZbEmW�H8(�Лd��*J��4�[�M�Y��~^FA)��v'!�,��ʠG���#�N=��\�y�40GlZI&7�fM�b��<)9��ğ,�~���n�ǓJ��(N���-�{���3��>�X]����~B�t����Kf@tWA�����s�Ӧ�0��fE iy�9�c}�H!�/�<Ԝq��M�ur��N�u���S�i� �B�Ka�{#�im�- �Dnnn���]ލƱ�5�n��Ⲃ���Ydyf*N����~���m�����71���7�1":����S�����!y���g�Β4I�]]O��������h3.MH���7���``���p���q{%v�}���C�����x��-����K~�8n��'��{{���B�Mחƿ�'�C'T��4'�f+���#.M{�z��HL~)���&-z��};\�Pa�0f{s̡^S�]�3�i�ܚ��=S����:�Ês�V��&ܧ0(6��A���5�m�b�!�ńM5k�l1��ݷr����죙?^՘F�. p=j���L��y��@���h`�%4WpPǒ�EDE�?��=�W�}�������@Zt�c3�t�3�ʸc�8�2+?�M8^���\3�ZC�!&�� �.�/wc�Ԙ�X�my1	�h��茀�Ff^b��5�~m���J���(��J�,�6��fΈ@��<�wr��7!122�͂[��N~t�}	a��͢eȦ���:v���+�qv4�
>Pp����ӳ�!ཌྷ~6��
�&NԻ}v�c|q�$�� �Ấk!xaO0�(B�E?pc�_?gx�λ�}pb�:~z������Q"�G��Eq�ݮ�����s����	+"����yڧ��x�w�C�E
4� |d��tR8��R2��b�MB�ˣ5K�Cg�S�ǢX,<NRs�y�kHH �_����iz^Ļ���LH[�)���!�1e��<���>{��Pq���>��M�i�(�e��s8�Э	a���x�Oͬ�tH�vbi�n+`2��'ʛb��@?�Yl~�\�N��l�iM�2��8o@�.�=�o��+�F8Z��+4�>����7��I�h-(�>ǃ�Ң`E�$B�����/)���2 �Z��*^� ���Zf`���P���1���ٍH��!i�IhA�/x�`��p��N��Y���~�Ў��Wen�o��~#hOҘ�m?�5�������><0��R��6���^��ʱ4��}+;~=�ߩ���M�W���(K��ݎ���U�e�+<�:�V+iF��d6ë�A�p��[� M,������@Ԅ��`���*g*Uײxvͥ5JT��
&�2��]@�8=X��Ц��A�;$���kY�����B���,V���� |VN��/�/r�G�Xʜ�֣���ᣠ|#a`ˁ�O���9i��@�&��ԧT<���A1D>i�-�:�>ؕQV�I�fxZfQ��h>��?��bx
Hj�D>'8����َ�5��%��]�s�^|�����"��p��u����:��}�v�������وJ�t�c�@�a�k��4��K�%"�l�02* ���K�AI�^�k�M��PL��2^���	�|R`X��`���i^�g� ���19X='���76�< ��9RF� ���{��^^�F�e��o-��_��xh��_�7�`f�gkV^s{��y��+�ى>61������kn����L��Md|�}+�!�g��;�&�{��)H �p�v�&`�����A4,��x��~d�mnӂ�*\�Dܺ;Wr2I�-� ���c`7��X�%�f�RrV=��&
������BP�������ae`T�:ܠ��Ŵ������6
������m��+}��@8L��������o���ll���@aHqёK�P O��|e><�L�����?�����8i�h�w���.��e�����0�� "�N5Z�ɏ 5�Iձ���$�C���մ�:n'���RU���
�ӟ�v`��y�������}BQ�m%>D�� ���8���_��rà<�*SO��b ˂M/��h�1�q{��>��<\�je���N��^I���wssl�:�3���IoߏG�%�N2�.9`db����vmO�\G
w��dZ��٫P��ЙU�6p"]|���~<��ld�
w(�'����K����E�Ȳ�v۳b�&���I^HJR����JJJX��55��H��Nk��m����2]>E2?�]BB¨���B�c,|����M�\�nnf��ot���$/YX4��$��\22����c�L|w�S�ϐ��o�����#�� �F^O"HFR��	bmN���'�����6�n|yPq���`1���BEur^K�(S[u��͛bI�|�;I�m5��%up��Ʈ�A�)S��'��X:t��׊������Rᕑ64�T�8��������{�F��n �[��G1Н�O�Z�|�ɯ%ʄoj�h�
�q��8�
���������UDn����]/��1mdDW>����˯	��%΍J�e]GKu!D$�v� ����n�΍(�ɕ���wxu�T��f��Jhk��^k��!�?$��H�����T^�.�S�J<���Y�����E��-G�!�ъ�{C�mhL�=
�d�1mj�)��~��~˿)
���R_TM���Fu���m���ڠ��UYv��kJ'>�_F���v��zW��ȟ�EFE5�z�9-��}+r�z��Y�/�n�V���Q�U��~�� ���t���LW ,��3V�.C�!l��K�9l�Ym���C;�;�Rm�k������7��>Q��6'NY�}��Y�Q�]���p�z�_RZ��r¿$��鵞cy;i��ӆm}"����u��3�6��ҋ����	���𤗕'��@J:T%U��:�JR�{�!Dċ`����W�w�뫙���c�=�K)�F1%OQ$� �*3�K��%���
��o���u��F�߷�t�w��5Q��6��n�����FlDAa��9�YMg�縥
H��ں:��G~?�W�:W�1]ߪxCj߾U�0�!Y�ui��Kk�Y~�d��׋�O���Mҫ�G���/��������`��-���ǐ��[XS�u�� @I�:����5�[���1�iU�5^��''U�Ǟ�\��ԎN�[��7+ೋ�-�߸%U'g��M���Ã�����fm��@���d���)vqo���m���`?w{/��Eժ��O��@
�m!���,��!┡��4�̗�������g�ȿk�.-)�$*;}��_m;RQ��|=� ��������ǎ$���v�^����؀ ,}��n#E�2\�t ��gQr	!u���Cg�|d7�*� q��jL$������-�ӓ�}:Gʌ�������&��(�}*ʰw�M��?x��J��f�/�ځ:~?��e�=T�{��6��:��+&v'��/���͇�M�o� ;�|��1�ݿ!T1�P�k��V9 ���'%���G��}�#��t���b��%�k*�s��rsY�fB�:$%��f?L��̚��#���4F��/\#�V��gG���ݙe33U��Y3�fst�E���W�o�kF%K�kFW�f���^@ڌ�N�����ˑ�b�7Cl ����
X��å�[U��h�~���hS�>�k�ۈ^��)��)�7ܟ5|!4��fS�����}�i��*5VTӨ��@�ٝ�"��˼q����q���BV8�w�L|sv1!N�籸�4��\�/��?��<���ƾ$ʖu�-![�Q)J��!Cd7#*[RJ�ɒ%{��/�KY��kvf��1~��y��y�����s�9˽\����}�?;̝�|u����'��'���'��k�ҳ,>
�l^EW��Ϳ�,������Q���t�2۟��) ��Rd��\i�,���/f��*�$<<���GN�Z���VO�I��ח���W���V��%)�.-����Wz��"���2G�䃨9�'�`���y�}B'+&�ƃ�?��.��hk��7�}��KZ��L�j��H���b>P���h���y����u)?"��i�	��vz���
������/t�Imɘ�l��Е<b�t���S��ޖ5����Ę���_KCp������ѯ;��ӓ�<�Д�q_^���>c��lӑ��ȢV���V�k)�U�̶�p)�t5COMU�^ʂ�:>b�Z������6�wj.�̬�p�w��مU c�_	��C��X����犿'2�tȢ�"�O�����$O�90a��]�]1�u��P���\�
�*���i��K��I($���ˤְ��zB����D������b��R[	�us�ߒ��~�NvJDIPuʴ�饞��oN�U0��>�Ut��)o��%�j�f���_ڥ�a�h+�!qw}6���,ǲ�x�s1���JLdu ��:}�����X�z �c ���b�ͮ����ܚ��H�y�]�'�S��7����[1p���GGG���ϝ�� B���s�����%y��4��`I*$|÷}p#���x� ת�˿iy:���	��-���� 	�����;�13�����T�=�K�����=,�U�d�ۅA	����8���s������?\�Nyd�@-�x�����R���ċ�J�Z("/Q�j>���h ���0¢A]�v� �� W����\g��)��=���ݟ^5�I���:�uyd=�]v0���D�8qw#�,.:}
ມ�t�w��>��t iR(1�Ë+�!� u�Ώ{�xd�&��������a��4�9'&�.{iɕL�E�h������ҳ��W�$[�S�-�����
K����}�;��FN�쏮�����F��k��=M��	' lV�^�2�3:1Qu�븙��T��x��T�zxkn^A���-2|�~G�Q��o�$���"���/_��;w�%�z�C��|XKSڗ�-�L�
�w�Iv���������>�H �����]s��ǔ�g������傿ezr���MK�X��O`i|ym�OU���\xJJJ�At�KI�_�qtr���"kv�k:���ɪ���3њ/�\�(>��:��aEC}�z�'-�yW����II1c���6�2D��hO��[j*�8����n��0��(~|��`xp���<���P��8�H�g�ɟp��)���&+܊F֪
�"q�������Uc��q��#��p�ZT���0��/s���;jLv��y�N�X���m���o=��i�����&������!����=R�l[4~��"W��"8�^�(��>�l��íyU}{�P*�y�3����L��Ê��_-±�1��@�o��Oy�:J&tv�`%�v�#��ɳ��(�ەi��H>�n�P���/�15c�v_�ȑOѵΓ`����u��B�^1:nld����lIjJA^�[zέ8��RJ'��cG�<ñz��[��c���/��W�q�kV'G�����
�y�����{��ܝ;���YS:�_6y�`�ړ�[����&�=�1M��Q�W�x�͖�O���O��^0A�����	r@l ��68�#����bk� O���Q���;�fCΪ��GW0%���{�?�z���QJ%���u���;"��_��}�O��٨8*���G����0�Jҳ��C���ѩ�W�������5�QvI7���a�B��9X\�U8����ޤ�����l��;��b�ep%X`�\l_eQ�ZY�Ћ��w��cs�P��?��7z����V��Z;��)v>���~��6���6��Omb�]�#�Y�����b��=��[a^�U޳n��q�E�u$Lbe�	925ݤW ����~u^�:�x�G� k��<*��IiD���8*'g���J��lt�[�輯���ˇߴc�0o_7_�VT<�W6ŰҤ
*7qm`*-�"�H��zŢ����.��C�~/���?��l �8A9�z�9zl�N|���}g�y��;Z����~����T��)�5����k5;I�S-�J�-Ku�|>	7�\~F\g[��L��4ӎ!T�q��ǵX ��&��F"1o��}���[E���c�?���M��TPs���tQo��I�>�W��#;ߨ��+���re+����b�ѳ��P_y�oـ"o�ҋX�S~���@�����^�0�x2�%�����&+h��U[��֐�o��2�E�Mq������ϟ�����NȺ�g�7
9�7a|��z���J:���Ј���a�-0�`eD���$*�yע�9�ߢ98\di[-9}��A-�o�M��[0q�j2(S3
4�����k��gP93�F�>K:��In��Ƥ��L�>(]兣TV�Q�lpI~��
/5K��B�ptB�3Vr�����m��/�8Q3C>bծe���Oܺ���De��j=��о�Ru��s;��v�+���ۭ�:�+8�}��0���D2+��QZ<�@��M���]�ˍ;J���*���Ė0�4�)��,NgA��M����4����y�۷�����9\����3AR���u�D�\ 8�*+b��(;�{�4p6�(V	��h��]m��j�-m��7��u�+Z��%�ˢ����ۧQ�'�+°,P��]�pOz�����4�9O�l��/) #?��1���d�dl��>��TW�~�HP�y<�a'<s뎕�8�9�3sSSS�x�Վ�\����QC
l�ڃ/�M ��	���p�L��{���u�0H�{�����4�y�N/l�ND��Wɷ�K���:,ך`l7ܦ�ޒî.֤WE��I`͇t�+)�>ü��@������e���e�^�x�Q8֛:*oJd�l1p�p�k���TFU�]	��[JE�߱{BgE�Σede��ɞV�L'�`ʳp
�^!ň�����3�RU( /R����}��(ۡ"���w�.ܟ��lǴ����������=C�ϟ?7��.�N�&��O��,Fi=� ����*��������S�uF��	(�瘓���O  ���m�6ǚb��#�����;�6v��M j�(�Q����@��e�.�C��iv��jb���p��'����ߥjٴϛ}����(��3tW��m����.I\���ݯm��ע�{F���U����̊�lG�@�vY�v�!Us���=$͡���NK�}��A7�&Mq�9{�ll�`ի��sƷ�WP��&���W���Y�w���x�����u <I��d�+�.�y�����+H����۳+%K��V~:����'�����p.yv��|�c굷��K�3���s�BW��W�yVU5a�b��+u�U�#ug��~ό1.0f�a��ʷ�G� ��J��������
aZٿ�}��
.�ui���0�
ܢ�;��3η�$O�ȧs �&;�m�Pq�2�~lt���T�Xԡ�]%�u�������+W��cc���wvE�&�یL����XJPvp^oyǷ�'��I�@_�2���Npɀt�4�=8�]�� 	J����W�`�n�Q��ο�����Xb�C��w�6e�v��3)�|:R�t[�f�Z���T�y��\�* ���j�ڷ�?�䷪4p�S�`^�t����m<�a��/��03//Ҝ���	�
��wl_�m}�����\�u!pf)n>d�n;���B��X-����	 ���5prJ��ԣ�4����CVx�CJC>���H��I�6n \���9]����	��(����v�̛��jH�G1��E,����U7溟��'��$p��۹��dѷ�ch8��.�_�]�lh[�<B��m{*Fm�p���)+3Sk�(�NN��h������ώj�`u4��K�7�W��C;7�%����0+��J�#����|,4.����h�P�po+�	�n��3"C��Oz5m�y�T�|����G���b7G�v�^��q=���Hy��~�W�ȣ	:^fq�<���A��3����">�_[[���C�y�M�c����E�m��6��B�q�պ�<�#<o������ۘ��]�_�n��	�"�|�����sk�A«���'��\�Pҍ8�+�{��з�dK�K��U� �Ȇ���FxZ��l��O��ﵡ��^�HX2MX8����7�L ]%�g HD���O�3�i��3�zd���F �
^�"����!EGk�c�j�g4�&&>��ྲ��r�g¹ׯ_��(��Up�?��Y�J��痷�y��d]H��II�0�}f��v*���uñ-VV���ɉ$�}>vP��j�[�Wϖ2�3��̃�����W�Ǽ�>�j���b2t�������d����^%��4�*wB�-ze�dj�7D��a���27r�^�.|t��k��`"�1�̜%N���W��)SL��Ρ��d��'�a���E��mx���򞤞ED��ҊN��9XAF���/n�p�:wD��\�N�n��r]�~�pؒ)�E}�C�R��e~��3��s(ע��V�V�`�� 	-v�+��0*��:fb� �h^�U�?��Y���:��������(.��9�n�H�n��J���);��@�ܻ�?����W?���K��)��;5�k-�ۗ�����qo0���%#�)��r���z��G�U�?�rX�5����<�8|:�޸�?~X㽘�qE��~mOȘ��o�n�7q2���i�������l�/4gw�!����[F?X�h�|��j�+Q�X��b�MTX�=h�����"^�٬J�
K�����RY�<�*��.�E�6�c�9���TĞ0��Oy�Bz|c���σop��Bt������ώØ�,���9���2��)3 �����u�
r,|xR����G���h�Ȣ;,b@D�om��^���eW��C�i���k��WCg0"��3^�.��ٰw۷�C��C��%�ɍ�l�"��T߯�����z�'S�x�L 5�SaZ�j��>�v��D`/����++-���|��=��x��e��ۂ3zF�~2��"zI��4�'�o�^H�!��P5�}:��̪ۙ}�cWMHT�yo��h_�h-�Tṫ�p)ы"�={D�qÙ�΁�s�	��N�f�.�%�z��*=n���o-.| FGw\��Xr�	8�6|)���P58�'ӗ��r�4���c}��$*��S&�{ok�;j7S�([ñɯu�j���P�� � ��5?۸]Ν����P�%�[���S��
��ث!�ÐK�Sf��w#��2�X0��=f����X;�?$�՚����|Ĩ�	���#�V�#�/����Y'�nM���yR� �5蛓ω�{�� ����ҁ�X�V��[��\�}�4q�d�u�h_��`]
�4�*�``
(s����/�}�?a�|�n����rW i���4�`�~xt�5��B�ԍQ�6m�������+�5�B\��]:����[p�2�X�|%CB��%��O�S8���`t��H)�+U��4��o���o�N� wW�i3;�S�O���L|s����wɬ��J�gJT�]7!�s�3'��	��GUr��y=�K�y�M�1�9���R��-=��4_E=[V�`4�AaF'�n�U��K���4����z����	}�BS��ޠ�>Z,�<[b}kM;�~}n{�������ϸ��������΍��Y�9Q�yE+N�	<���I�'6=W����Nʄ�CU%��LhrC�6j9fj��m.�JY"<�a3�IEK����`��4��r�P4�b�A���]�L�p'�0o//;p���n:�/1rHD��uFcb[���&�� $(�UMj�eBOV��L���B�S�_y�S�!��p1�(8>����	���S�������;-�_b@���Oj
�%�����Sk(��y���Z5R-�5�z��ǉ�ffAǷUx�@0swX�����#�Jt��
�����9AH�j"wb��$'C�em�?��y�B��xV��*J��q����#5WZ� ��(�t>M��Х�I!b�qu�W�����I����a`C�Q��M�f����y)��@ϩ�R<�qA�Αh����@�)ɍ�h;�SN��$QQQ��m�:�8Q		D�+��3!�1�=����5�Մ����9����Sw# "�����˄�2��r�H���=9?sCK;�*M*���"�]�Ռ���L��DQ���&U�օV&4 nA�;�o8I����0�ާTK���z+�cd ���v�$f

\3�����DNI�����S�"��-r�T��3*
vUw���U�k�e%�h����5n�Iw=�_V������L�V�	̼Cɇ���E���[8����|�svv|����w���}�M��OKܯY4&�9�d�>He�ɫ�z�!D�3C�4PC*Kj���M�����Y��B�@��2�zդf�@�v�A`�z��� i��5�4�!�=2ݎ�[��!��.�JW��[J���zX5�8���6	�=�>s�_^Ƅ,�	���)I�V}��`>�-�>V	բ"�R	���rB`-R+���V��h���h.����1Z����h潁Nk?\);�>N�e�������hhh�k�Iiw��a��Z��2�QeW������:L?��GH.Q5+dD=�н@x¨��������{K��B-�t�m�%'�U�,v���Nq��LjnJNt���l�XZ�c�K������#�q�la���CĐ�"��]%�)�"��8��?2g����2������U.�����[�ۈ���}*7,4n��>X��Q��T&J�<�≷M'z����!�X�kV����7�����H��:�(���l�Ok�a�����A��Z��m/(Q�S�;����;���;&r׵A7�%�/��:{�-~q��}\�a�P���0Ne�GV�h��+�O�|��\[U99��V��y�#}0/ަ�ˍ2u¹�#!M3Β
��y��\*��Jk6��y�����?	��	u<�oEԢN�Η��_j��O#�b������)�Dp>W����?����v�����
(z�)���1����� �����.ww��h"�YVzv�4��גKZ<�0�M�ԏMm����ۜ:��f l\X���DU��1Ohh\����>���4�w��>�!�7��������r�5�.������@�;<x 7����M/r�9�<�!�<�HS[r����)/��{�)�66��/-����*��a��L ��yM��%����a
�a�x[V��DA"���YVr��he�:�ŝw�'�=a��ݎ��W�OZ��!}���?�o�ܟ���H��Hi���/{���s���B��y����c�F����K�9�U��QAA�U�l@5RaP���� �j� �w�r�n��@��P�C�\��^��f��C��.�*�S�Z �=	*"�f1��Ǐ`X���h�~�\�?�%ka��C����I�I[�>�|�z{����3f�
�ߍ/ǡ��@�p.�)��V��d�b>s�=sQ����~�*wrUT�`QH��2ͯt��x���}���-u[K������J����ޫ�0W2/O_��?��)e5s���%�,�]=�=�L͛���~�2σK��_ޭ߿ך��ՙ��� �k�Q�`1O�V��^����?(�۳��_䂣��0�O3�`�8'�T���@(�6frr�	���"A�`�=��g<	p���\:9Pc�B[Z�}�({#cEԀ�N�bҡ7�P��,��/i�����7���L�oN�����5
mAXٹ�9��C���J��ր��M���]G,={���͇��W#fp����P[���_]1��Zfvvj�wt�ԲM�����e}��Ɵe�}�����}��VȌ\���bk�O=xL�	�mV��6�+(�H$��[�u�=����A=K܇�a����.�$7�e^�����_���4�{�,p.��}�i^��S�x}M���}�����J��6�U���{�{-�s�cY�����o�T�4����k�wD����:�N����1�LTn�V��7� �&cB�����7�:,\ ���=ѣ��o�CrC�`�S'�0��͜h�2��]��Ӓ�����]$��z(%��¯rk��,�%����('���Ǫ|$×��B��펄�e�5���'&c�͢*����a�'0������2���@a���0�?��6�$���I��AФj�f���=��Ɲ4Y���� ��:�P���D��AH������k/i����-~�{����ճ(uNf�<�+l>X-�-j�"2c�k�m:�q^?���di��S���g&j�l�څ��PjLb�.����K���]�Xk��<���0���D������U�K�+�?�5�	Pf���NŨ9�_fV�da�Wy�V��\ �T���Q��в�|���c�-��/0���0�۷U�XyO.��k�F!����r���*wV�V[ه�D��m-͙�:W��+ѩ���8��'�ç�G��DA�Q���f``����>������4�=��ƌ���<�3^��q��Z��:L�UD�u-eW?Մ���w��FK=�g�>�J��Ӻ���%S��v�/��U�����\�jG�;�%���c�\�ٸ�=�iZ��灠��	�v�����'��a��N��!�Xcx�Mm�Kgo�k�'&0�'@,1]��R5����e��|dg���C���N'T�WX�%�g,2��gk������sg�#K��-��Z�V���B����=RF��>9h�8�*{'���Z@���mD��n>"�@�D�r�5�偐h������i.��������~�̔�C��'�8:����QK�n)x�_K������Hœ��O��k
{z������?i��\o���4�ٱe��Q__�/��X�!�(s������2��zFTH��1z�z�vU�e�}e��S��'*����&֨ݳ��'C�ڡ��psCSgydHj������Ѡܝ�w��OU�k�t�Ί0p�{F�ܘ�Ep1����m��^)�`\���'��lM���0�}4�+·���+w*����*;s��Y&ם�ǗX��Ĕ����D�<��+Q.��B͓�����wb�թ�
$�v �B�y^��3+v������6[�}g�>5uo퐌�Ɨ��E��#�����/��o)�v���/���"+�V��WN�3��.�	}�|�X�/k�s�'Z~����Z!,�d�C꧈� ���ܲ������٢t������AJ�˗�:I*��D���b����̴�ƌڸׯ���$~�Bq\���B�qqF���C!���*�Ŭ����3��^B2��@6<���@�$s~�����[�����[�Y)�j��7������<VG�V��SflC'0jP��\� �0�-���yW)��B�BI�p:�d@���(�OL;�qޏn��] /�^me�$5-M�s^��Ųi��u�S����̳�aH��Q��͂����vvv��ȸ}�)��$��������X)k]��	�V^Tr���ܻ�ec�nAֿZP1���f�_�X:?�lv-C;�<��?�Q@+�h�%v^Xx�÷Yϱ�QSuZ�X����h3}�߁�QHۧ ���׬g��T�y���~��^�~���1��EeZDFtl�\�(�Bx�@"K�a$���d����Q#��1��!��Ã�ܱ�����$?��{m�lcd���O��P��9�%�/�سb��{�	'(Wi�/�>ػh{�B�hå���35�)�É��!:�F��{zz���k~�uW��J �E_��K��d|��C��Y���f�d�� �D�f�lh<��s&A}���e�g�/`�)т/;�/50�0opJ\�7��M�a��<�6Ã�v���b�I*�q<��g٤#Iu!�k��eJs��9A�;�``�to{��K*8So���D�O������&YZ�5p.���+b��Sz|��T�S�����Z���*ޅ�[���r������no�gu�0C���o��y5ҩk۬��d"^��Oz���Wc��ZTb��x[m�7Q~�e�2��4O���p��f���.�����v�,cR���S�Z�vLe��2�}�A�Q�I��Kb�����+83�� **���q�Y�Y��L8�Ï�g;/̾�W�cd���]V*�)���"�jJp_\��#��|�hU�+���B}/��k��rw�jg"ۼA���T��Qۖ�}�	���4'�� ��b�Q�=
��Y����x�� ������]�Ir��O�#eџ��_a���_v~��Ѫ��������g�Bz�DK�(mX�y"����Y��ƥC�ޅ���q��`����ޛ>���Q�kѠ�I��sl�nO�4��R���Ë�����\:w���f�$�@߭�Or��{��)�L�l�lB��^1�@�:̪8*�+w�霫3��+�kf�G�b�������F�-�P6"��~?��˗/��iq⢎�
�����
`��H~1*���s�c~k���_B8�_��5�P�t�
n?%�>��y|�ǒw��)5�����U�YGNR&����E���ơy�]{�ȱ/���}�rq�!�v�*����@��Y9@M�ׄY���� �i;���o���'6�aQ{E������.o��Og>���y�׿4����(���ڗ�
�,��1�X�k�2�p�W�TM'�,��=߱Vf���Y���&gkF:2���8�����ozF�.��� �ϫ`��ӹ�5Ҳ���t}Tԇ�%�tO��o1,"�Q���˖��3���!D���)w�<걓!~u��,E�M��&��̓�������������j�***z8R�ֽs��,S�&�Zk^t3�oA|צ���Ԛ�5�m�Q�X:u�:L�3�@��	O%�TvnLu�#��� ���mu!N2���c☶��w��a$����	�J<v[%��8��x���]����3�s�#(�5�hJ�����I�C*J]j'R��)�<�wt�bT_I5L�X��{�ߋ��+�����[Iٶ:Zi�߰�$Y�J��ɽ��Q&2?٣�ni{���Y�Ł�D��ۦ�!�v��̐��pcH�
�%Oz�Fw�:J�8I�.���4������Qa̱��QC�Sz��mc���Y�?��ٷ��C�X���j¥Q�'��İ>�-Τ��&��/�<gD�!�S6t`n�{�f$�B�k0�j�v}�S�\,�%�ֹ���0%����(]t��}�^`�����aѓMM��萫_�<6m�=�R�p��/�'+)����v�QbxV:�h���xڹţ��UO �FA��B1��>����9��ӗ�IT�bz�?����K�hH�9���0ٸ���g0 x�` N����;�K�'�6�BS��}A�������&rʙ*�������0�����5��*m�A�����i�)��/���*����U���!
�%ۑ]�E�w�?7${Pw���Մ��� {K�0�|�-�wݷ!�Y�}nw����D�{x�RHp��7X@l{Qwj�+��pq�K���-���ѧy��c���Py���۾�׀~X�W�1� �t�o�e`��������HhK�a`A��~+G�&+�s{��5�l:ȅ��(��",ly�u�����k�Aq,Ӆ��9H�'ԝ�xwS_�K�&�����ˇ?����lcx+\aA��«��A*�N����v�XVy���	�@"?��*����M�t�:��1�BCu�o.@��l�S�L\g�5ts!{��zͮ�.��Naf�l)T�58��	�q�0w�x�Y�NŹQ|FY���<8�Y���Y�����;��������(���u^Cu?-ɢ��@Xx������h�'��h��j]#�=�ìAG��ru��1�M�w��i֐� P�|�&V��� �e�V/8�Q���Q2�Q����� � �c]�i�[bw�<�$�"�i>D�uf0W]I��喭pY�c�s-�d�o����A��vr�պ
�����:�d��I���!�x���ݲD�z5����ŁȌE&���g�sP8�:���������"A#�e3&g��� �7�%;�$sw��	;R��[���]Y���X����W��JϺo��I�������
������E.��!���Q����i##w?[�|�y�9	�O��*J���#^3�/��R����� �|m�k)N��UO���N�b�S_����(T��D������b�,^�Ws����i��&� o�1=7����_AԌ��Cܧ�N	�z��n��G��e-M��4�)~�Io��/�ggg9�N�3L�6C�sr$l�뚘	�"E����Y�[b7E[�>!K.l<^(�S��o�X�W|�`o������c9�|9�C>����Dm\tb�}���� "o����M�M�jM0�'h�@$���}3FD/��G���Vh�r�f��)��R������<���!�Џ߱]/$���N�r��u��i�'.�}��8م�Z�ǔӛ�oŋ����u�\��pttt�c�s\a��C��Ի�]ɩS-*�c_���'�� ��7��"p���P��d���F�P���@�� ��^���3y�-�������lUB�`��O�,�]��$6�o�{�,F&��f\_����� ���v5�������+�,95
�<��:s�&r�ٳ�ᤀ��)�~,���d���)y�)���[v
l2=����i��������nx� � ��1?�ف��G)K��NR�Ic�"'��و�8��������@����0\�&ɞ�S�a9�'4*�@Z��G�ZS�!s�XJ���W̾��KO��I�<���
��~���֩�
=���ߍ\���4�qׂK`�K
��𼢥I���w�c�\�W&���n��̗�V0��T��5��3|�8��x 2D $?1��R��yK7��U�;A��n����S�/^�K�'�t�J'iW
�z�9?�e�]��h����燅jr?\.�4�LY��;K⳺KB޺q�؆��CsZ00d�ќ����/+�����G���c���7�پ~Z݅�I<�L�@�ƣ|�D#��2]5��x���.�)�zk�-�z�68][��7~�4���I�( ��!�4|j�F� �1l^}R��� C ��5��ߐ8�^jD�jii�U�uO�^f���r�u�� v-�q�9��cD����J/�%�)����M�=����X�f'�JcH������6��ZXٔ;�Z�	�?�Å�d��p�杤���o���B��M�-rn�ފ`$�R'����Q�8̿f�귝�����;��~�e}�{�чe���@�[����3~hӟI����
w��-��rU�;��T}߀�|�.R 5�0k��q���̥gu)���ך8�=F��kIה _�	�/r�+|6һ��j��i�]�D�L�<��6NU�M��Czz4�<<.Vo�Y��}�����Λ�'&?����
�h���.�>+��#��X���v�������ѭ��Q��Ar�߄hc#.�^�&��:Q���빹Il�PhF���TJ+[M��Bۖ�G�/v��o�~�3�kH�soh S�𬬬 2ڮ.&����8����/�qr:�|D:ɘ�.���B�#�	A_Ȣ$P���V�|�2$lB����߿�f_9���t4�������Ս�� �R��PFTWUS�`�bQ���R[�|*%�+j�AJ�i��R?9�V�	��T;0c'Z���h�k����O�=e;�� ax�0�|��Zס��L�����>�%@����b�R���!�y�pN�Ć�s�^��&UZ�W���:�G�G	ø�`Z�W�6�4G�S���} l����l��������e~Ḡ���
�����
ѱ�E�)&��"/����� T8���:C4��'C8��cT(�w��ѵ4��`vR�qug?ec|���΄�YCݎ�1��@���9-|��o��� �s'4���s�f�VH(_>��M���ؤ��C} BS�]j�J.(88\A��3�ɴrgMt��[}�<�7���>�����ş���o.L�M����ZY l,+���y����+���P�����w�4���r��hp"�"Z!]�}F�$��/2�T_ �Jqċ��W��՚���rzsZ�hÏz�GY���� �N��|��T�&����`���<j*k�.[t_ap?�܅�ՠM"2i3˾l�'�.�Rl!滬�O�jv�*���i���KJJJ������C|����k��#"I�1 �3_1�@֓D��zB�Ł��V��ꓚr��I�dA݁��'0��G,�y:�U|��'lT8�'Ʝ��� ��/s����a0$={�bO����i��Snaz��<h�x54r��K��>g421є�o���T0�WtOW#j�33[�~� �K��{��*?/�����3�M2�Τ�'`���k�1�5a�,@���]���$�c� �1�5��QJ��4�o���`�	!��Q�J���U-��By�� �퍒Gh)^�R�����{�'!��(�$�Љ@�zL"x�~�L��$~\=g�y�J=�wI���n%�X
0"�P̣�4ّ|5䜊������5�2^�2<xw��`�|�Z�����(�x��Қ�~{�B>v��b��}D������֚gE�j7o@E��z��r@�*c��E�|�*·L1�e���M ��;���A�@�x��)���1�IlpЙ�P��'z�9I6�(B���W��Mm�O���<
?{� 'sѷ:=���Up�|��^����R���j�3����5�Q;wt/q�f�@��}WO�z��B�e*���J�!xAF u �s�\�΀H:�z�W�2dKW�07�bZ��M���&����i�ϥ���8�a����Z,�`���[�m'-55N��ϟ����kU1V>��+���|��w%��K�['��1��d��7��<xнC�)��/^�l����`3��ݿ�j+��Q�&5�@/��u�%�0**Oh�HNh4��/&��8��EҀ�Q�Ph��.����P�@~Ũx��	/hK�G�y�F�D�~&*�1�]�C�V�̌]>��t��}���'�M_җ^$�k?b �+��G��;�A�a��F����տ���ex�h���p)�r�G{���(=��ʯ�@�S���߁�2�������2���dt��P�ݒG@�m�9�˾2�Tm�$c�^Ȉ2�[�k~D��-���EN���� �gk9��sWa��p�Xo�	n_J^=&��|!�}��NZ��w��x�I���@H������?:���w{��vP��٢xͧ��y3JK�\���e�YۭK�kN �[]��q�~�n
;
24WDt
F���l�I�UT���X��_��`�1����^DLfx.q�L����ά�.���w%&`�ϒ
z!��?;9P�.L��&g�f%6��x���;7��EHwku��ʰ���3�rc#9�}�y�7HC�@�\�<��+�����37�>��P��h{�	�ZJb�ˑQ<ƭ��=�}�a'��7`�& �<ԅ��{���ׯC<���#�y;�_�Ek�'O�`�Ǚ�����v�F�˓$9竒�g/�o1lQ���bu�K�$�,�����g��
����u5��m?����}PTB$���e����4���Ō�r%<�@�?U���ll���"�S�׮�@��֢k�
R5���S���_y��ܪ������1 8Z�<����b�O��r���4�m0�����L	��/���pSB*?�T�'W�=��m��L�)�<��/ ���l#u�~i�x��F3�N&�@�[�E�Y���'����	����m0a�X���zlZ�3��/;�i��{���G.��T�?Ow?���"��K�3�-Nť���	P�|cܳqś��Cۏ�����{G���p����l� �{���B���/\G)�0E��Q�����ua5�/,*)!qA�ĥhW�+}N���Җ�}���W�.OdP��W>�u�r���;�eQ$3B��9YT�ej���Dz���Ң1Rj�{�.��7Ѝ�h��E�3Q����*�E����:,`@A�RwT�Tϱ�����
�����Ձ@��h��������dL0O��޼y#e����I~����d6^�,#��� ���
���X��[�gK��;^�(d�|���,�@?�vb��N�������U�6}=q��������kǫx�,�������ߪ�J1!��t[1�Cc^?�u���Ԕݼ*�P��/�K���l^J�1�lcGj��Ph��s�%!�I��f#���&$j�'_��0�� ��aLq ڵ.�>>>lllv*-s�hbp���.�����:��]��"�N��=��>Hf��d�L�yy
и��W*��I�	���W-�m|Jw-�qJ�x�,�t��=O4`k�;&�� I|�{�F2�1M�#�(d�������r��'���jQ	��L4��>�p����1|C@�,�޽{g񛼿�P�3�R�b{}��cZ�Z>ǏQ��"�tmθl�pH�m���i=� �̌�s�x!պ���,=(��������������vk�����H8��o{��ګ@x�n�����/ϿRh����/�r�F���p�$_�k{;@4��B�o#��ң�^���M�_��B/��d��(�u���Ƀφ���`e�:�wW�A�l�t�E�Z �c%1�o[�?�_�?~�w�C��!�Z=�54V�W�*ce��p�Y��w�벲@�cw�x�F����DJk�}S<O.��d^�^��6�Y<&� �@#1
�q��u���l"|�__���T���y �{�?���$1JH�QD����I*I)	W�dK�mF-�B�)KD�fߕ�e,ٷ����`�������|~�fy���<�}��߯s�c��E5��s�����4�:�k����^a4����zT`o��F�Қ?g"
Z�s�������Uh�Մj�s\�?P��	"���S0Ƕ�D���m�y1`���>�F��~l�l@4t���ׯ�r�ee��}HM���C;~��iof���y�}�{���jCt��d��f������p�f�o:�ε���:)�ѯI�����)��F��˗������byn8��7�?�x�<]]�e���vF�w�� Ȯ2�%k�ѸC�L(\���i���_U=�[ꍢ��i�3���E.?{>�L�͕��WUW'�G��kN�QO� �J�M�=�c��?�Q�
b��.�)D�*e��}0im�뭲�^�ݻ��
�mVf�]t�	{�C�T6=�#��b�m�@��8�y}#.\J�(������tZ��8�}ԡ�c��z���ֻ�]Yg���9^�+�ԕG�������1�e�Q�+uQu�n�[���ԃh)L��TQ����BC�IRG�dkS���}8�)���/��|���VK�F�}�M���?~�I�y���j���<���%�Ç-SvI�U/y�0⊊T;�tpo07�H_ڷ����}>��u����;��JDg�zp���\>>8��	�1�2����C�2F��y��.}Ա�����`�*��U��V�IG(���7�،H$��y���5핽�{v-��V8��#��y�?O��C�ﳂ���fqd�?O�O~�J�Vݜ٧�j\�C��C���(C�D�ÁW11�gz��7����r7�̏��	k̻}�vs�%a�1J����r�I~Ӽ���G�p��//d㐿�a�]-(ɥ��8W�ʂ�]<ꀝ��Ht���9���@�2�W��Ӗ��R�y�������7Ou�5�\:M�3�z�&���δ8���[r���m�G�:�+�|s�S��B�1�̤����X&R�a�l���c]K���߿_��\~m�x�p[C������Mt�/R��ƹ���{�Jᗍ���	�'��rᲹ�]`lB����Ab]�t��[��f<���\i�X���T�b������x�|��Z���K�v� RyF\�3�_;� U[��WO�i�n���s~��]�l[f��}���Z�3�O3�5�"W��LL��@���猡U�ʤn�pĉ�v,��J~���hV�,�n�%�wu	 }�c ���u˘DV�_�}NI!�������E_���šw~�����ae)�K�$b���ͮ����.��CQ�٬#O6�W�w�85v
�.抷��V�}�7� ]�Rϵ$p�fr���گ,�������E�<��_�m�<r�-'IIH�RX��0��Qn���92�� I?|��fs�,�7ױ�������y�Č����(��y��^XʩV������hd��C����N���˘���;\��̴��KJJjal��O��p;''DZzQ�-s.h�_l��A�u����oHAe�� ��F�B�E�+p���1v��*$'hjùA�����$'&~eCE+�g�Z<)�Z4M�d�}oG���k�/�F�����k�9��/�pXg.���{���|��{�Ƀ�A�x�Y�)Ni*�h6�@�q|�ũs�5���.�'q��	�Xq���mIz�����f�Nߕ~k;^QQ9�r���V)D��G��� ���3	�K ��cU�-�Gxz�}du)g�H�t?"�U�70x���gKm��m3���=���ɕu��/!2X���($��)84����)�����e`U������4�Ik���ho&F���d
D��0gA�R�fx�A|ڈ����Q*����B�EWUU�577�X|��xt�=-�No�>�s���5k���P�:aBԗWϛ����ͨ�q�w|���nD�8v,9��]N�,{��-F{s�5-��x�YHȗ>�r��ƚ�]�zY�����*���E��s�_�� e�L��|����{����=UVRR
1���m��vv.��r9�U��*E��Fq�
%_��qbĨ����V��ҠF)n��D�����ׁ�t�Cᡠ���үgŷ$v�ڴ\t�y��qat۔{x���<r����3�T�' ���M3�Z�غQNE�$n��/pPN1�v=(X�����ɹ�<��줓�pK�8&x��/. ��垹�K��)�d��h}����t���	+��ay^e��x��y;�$Ҏo���uh�{���.�y�����,7\�L.i�"��}d|5��dg~� ]�;ꃑ�sĮ,�	Ц�\��m�v�'�,L�!B>92rN�ڕ+�E}�eCb5��ʒn�Wi�7�EG�M�'~A��+���'prtjuu���V����{�����iD�k;�r�,e�  � ��6T���!.��#s����@��fo⽫_8�U�q>4���a��k�/r�=��zv�e(�M����y�'7Z�͉X`c�^�/��j��&6K���g��� 6��M*9οE�n{�U9��Ӹ;TVa��*6@�����V�Nc	��*B�`v�8R�tM^R&D�xqb�����m"��䩺h�+Spʫkm��;2y��m��L�Z��?�e�Y�����Y�c��l�N�42�p�^ �)m�����	��'?�V�S,��kR=Fmh#�T^���c�i
���(�R5�-M��C���=$�5fu^xb�0��<�+���V���"dC ��z�P���P�0V��M!���Rv&K��ϗ�h0���#���^�:�j�	�C����gS��3~(E�8�P��RgO.*]~�YZ�t��N�G/ҷ&WrӜB���a��`��zn_p���R�D�#���8:�<�)��\<�6���R�;�:vM���x>R3D�����~wik?���s�g�����~n�]CY�`p�0�Y�Q�^���K= e1 6�P�FX(d$n�W,�vޏ���bw���5��f���=KT?N[�9C"4�+�#Ԇ��c5B��fLcp��ㆀ�;P���R�t\U�X!v�b���j�(k��5^6D��D���<����gz+h6��~ h�Z�Ї�Wf�.�k�X�;����{���M��&������g�JB})J�ugs�;��a;@�N:�.x4n��iCZGHA@���#�g�7��9Ϲ��vRx	C[J3be�J�D���0�q��
\��C)y�B��rӀ������}g�hd�� TNrNB3k�z>�o\o3w[L�0�K����7�NX+��OI>`��QuI����_���}G��gϞ%�#�h��`?��C��d	;O�pa��Ʒ��&!��Gx-�YI:k�Y%���j8��w2~WC;�6�>yH,�dti�3A�}q�ͱ��z��L�6���G8��~zn�1�-_˄\��L��c������XG���˲�ӗ�~�{ �/���	�� U���#�-
���܈)L��U�	kN�\G����*���)�ޮƕ_���0���xi��K���B�7�kMoL�i�MW�G��f����h�ꡕA,�u��jc�k�8�x�i��mƄ|ּ����9�����n2G�XSSӷ<��Pp��%
\Bʍ�CMn�8�����q��^�KT��ɴ��!l��
Sީ������y�2�R�����
¯�ѝ�̓wV� ���*������ͮ�i0D>������}�b�LK�Ӿu=X�W�jR�c4�5�MtBC�۵��*�y������������2G��1b*�3�\'� Y+�1�{�&�"��th�(Dw���� ����&	Ʃ��6���b2<��M�«�������� �Ѓ�s������+Aw���,6�B��JK?�*eg��,�X���~��̣��	�7�E8�<yy��i���-'M�`�6B�Og������P�����<k��� �H��sͷ�~���(J4�Nކ�hiɽ=q�m�K�q�E�BM�ݩ�c�=~U�����"�k�k�`�Y�P?|��ѭ#����w�@�O�^o����2*�٣������C�{�mǂ�F�`_C���΅�A�Q�oQ��n|Lr���-=M*)Q�
O��G�͡��S��^ma�N�<��U~-Mie�ز��/��h�*�r�'5Z_>^��J��Z�"�
� �Y՛lKƥq�1䎴:�o�Ru�_8ć��w��}��b����[Y)A�o�c%���z�N�p}M]��";���5�i��1A�$��6ё.���$=���в���S�N����z6�O����@���K۹�?tu]��mV�"���_�� ������6�j�]nĕEv����%ie��8�"��3�k�A�/�xi
+�5��W�=�~�޸�C�Q,C��G�� gY��A r]πN,�{D�)~f���n�ȟ2P[>�	�+b���E��� s�̺)FW���{Ij�~y�g/�g�u��X;p�������z���|Y�cدך�c�R�����]�B��a�������$ء���,����ϝ]
,�Z,q��\q3	z0�x!����7���Z0m��d��n-�F�[��)�9�7�JI�{v�<��C�,P���s�U�6��q�D�w���.O߷�?]�؎�n�����(Q��O����,��	��p,�,_��*Z_c������o������\X�uX����GBG�����5$��`w��U�[Y/d	;K�9�p1ye��DkR��x���-�0��ck�4�?�; n.�A\��[�m����WL��TQ�TI�퍲��lb/(dM�����ҕAn-��d�93����n��*�}��^x���ܻ#瘗x�9�fv�\���	+���9טI������=���D��aYJ�b�B�z��-6�.ԃ>�P$W�b�ʢh	5���$�Fx���,���{��}�T��EF���Њ1�C�1��|���*�7��A�8�61�=�F�]&�]sH����L����U�kfJ=�� dK�s��x����;r>��7-�O�(��H)m�z��c�	Y��7�F.��U��s��yU�P6PH<Ȍ��r0�l�J�� ԛ�i�"��y$y�����Ҳ'Ь�e�y=K��<�;o7g3ؘ�OgGGQMuk{;l3}Ķ��9�k��3�X�-u�=���.��Y5��m�e?�f�,-�+�<�!�k'�&�R-?`7�uR�=��8�xM�g୺���g3��N[��Q._O�@�{�����&���MО[$*��,7�����-�-j�Zxz=>!��bf�M7 �yƠ�� $��'#]�g@�>�*����+ES�QF�Sj�w�	 Ge����"��;��)�ƴ=>Al�êշ,�Y���M�m���C���g�@��h�!�.�#����.w���v?ڌ��N�07ڊ&��48K�<��Џ��H�M�$݀��b�21QQ6~{��'��`E���&���y��J��2�5z��\w�G��_�.Vd��U�?L���Ҟ�<�pδWO%&��SX��~֚���t�B��0<I�~B)BsAĞɁ�������J��g3��U �:��2�ĥ?~���Sa�ɕ�1.01v�	���+�g��Z$�Յ�r&왹8�3���Y�5Rƫ뱧ao6�n���D	И0�E@��:�s�O�˳�������_ ����2k����K1�H��L�B|*�3����MN���)�Z�
�!�On-F���ZV1,Tg
��I�a�*�������g��a�XbCE�Z_��8x���k�}��^!$M=jB��X>�y�;�����c��*Qv»�,�(7܆��r�T���}���2QL�خ���JղC4��L��Օ:@�iBl��ҽ��f�G��n�w'	g��~ ��H�pl�]�>�}ǡ
�7�-,�7c8;����A����"U2����t5G������V֖���QT��g+o��]V�M-�;�ş���`dW��0S�)80�_�B ��Ff`����NW`��{̂R׳�%�QZewz��b�7!z��8X\�O���t�17.�C��/u�����1�u|��8f���}8��f�`�=�p2������2�����e_�m@
�z�K�����2	O���>��R��<�pہ���ivp����ո��O����	��f��Ԙ$(5`�m��v������+��~����F�|u3�����DkRH���Q�����}���g���.v�w��Q'E�0����=WZ�b�ٷ��?�/K@�y�}"���5 I�q��r��G����M[e���܉if�(�S���\(���JuC�o���vr� @GXz�|�Tt½:��mQ�����4ȡl9�~Jе�s8�<����8l��%�ǉ�Yi��.����8����Z@�q��z3�P�������(j��^	B�آ)��\���Yk���j\-��T1��Qz��~f�(p�͎0����}Lj�;K��7ޚi�,�.զ����B�56.*�*P�����'���I�;��m�࿷I�A�qޭV�Jd�����Ώi�Y���a��a�b9�X��X���|NL��D���"�"0�(�Sw��	轑��k;��^r��d����9�����m}�S�Ѝ��N��$i/�]��c��9B?����P���E�k��9�CI��
���
����������hJe\���%p���nd��KV�mf��.�hJI����G��?��(9`l`?4��F�|��s���7���z!Z�	��dC�����jO��!*Pfs�Tmu��z�N����j�����`�������I�3����Y�*Zs��������kI�Vȵj�H<�����=�߳&�V�{��Amhl-D�%a���K�Z����*_��m`����?�Ў��C�{� 6��	�^ha�r\��_�oi��9�ss_��� ]��in�1�*������͜���1�(�þ��`�ֱ%c�APel�;���`��*X�톖\nR�4��B[�~�@>�rK�ݮ?�UY��(�F����E�p1��f�!q^��z]��S�=}�4˧�|��8�2�U��Wvu ���\&4[-��-��3�� �W���V���A��ak�q�?�[-����yo��9�w�X�����3��Z��ʀw�S�}޹�**	�+dC�;|�W2�PhFp�B��b����#>�,�T�>�3mR�.�dզd�'�6�'>���L{�nĴح�2
�Y�&#���NC���:4Ó�<v��&Zyц�L{Kh?��J5�Vw�>?�7�˃��\����ݞ��S�l�컞��!
�ct��^��c4���{�|߾!�
�$e�s�5X�3���k�&6�y/���˘���m����R5��i'�'$�lT}8�s:��Y�JV-��5�-�;'2���텗p��o�"��s�1J�@���E���B���b���.�.��氓�����o�03ޏy�6�p1	T6����""���Z��ݯG�g�졕�e�+�۷%���]:��qSz�K�z)�	�'MhyIN�Cֵ�t*�gk�z������'�����t��s �Z���D+
\�>c�Mb��:t�E���<(�������]�/%J� =��;����/���!Ͼ�c|���]�S���o�ɍQ�?>\���@����a.�K�Կ{}�6td��S�c�w�lWR�}ѐ���5nD��)�n�@f@l��,��Sg��he�4�g��\�ڢ�yC:=m��`�nK��ƺT���!W����l�W�C�Sto��ʚ7�_�2����O��9�E�1�M���������3��٩v;ҩp���Ii�����6�1�{�EwfY���H�� >�u*�}�
[-G�'^�U��R��!v�!�VwW��U��*����51N#�,��G��fP8�XB]��i���ʵ�G��f�����[r��'H�[z,�W ��OT� !I;RE;2�`y��R��XʉG����Y9��ӡk�Pf���܍6J�o�r�JF��8j���o�h�^���W���4�d	�4�����wy���ȱ*=	��'��䋱�6Q$�<"�&ڒ}�V������g�V�G����	fq�x_�ð��
���?_ڹ�o©WoY���q(�z�F��:$�˿���HP��}�Y�����A/g��*�z���4�;��ӭ ����@���i_��Y��NW�,�������<��� �� �^M��+��=y���VW��:�35K��}-�����7��.`ֳo��I��ȧ���:�J�*�R�����Klp���2@�}�
�M�*�ӷ\�.ڛ�>_+�B�9M�mc��aq.�J"u�G}��Q�>��C�9���7�xtn�����:8�_l�A��~û�����
��h�2)���N�x3�p-G�>Yлx�;DF������^{��ǍϮ'Y�ב�N�܌�c�:���^�v~��Dk��E����~��� �;P��7�R������������/r���T��H����R�j�mO�������D�-�[)R���,Zv^�x�� /�1���D����Q_*p�@�2H���ojZ�;�) w��T�{�B ��|}�3�vݮ��	hއ�C���B>�TV����D*��m�p�ҾmP])e�YM_�X�{ǾS�&lU�G��Q==44G�~0���J�p�p�mt*��RJc��Ix~Ơ���8!�O,���4�}��!i���������%Z.�s�o	
T$�8�Y}�P�f���,��!�}�:��<=��~��,bawEnա"-[�U,r���^.)Q/�Z:�����~Pr��tqҝ�g��`2{��}A�e����2;���<�8Ű��}:��g� TD?\��wW�+�U<4� �tR�![�~�ںm�!����8�mی3_���:qsź�ë��no/��[0���=�=o�e1�m��AQ�=^�V���1-�Q�K!���K���{�H=������ U��S
�S�u�����:�Q�xk���_�-c�q�A���G���w9n��$����B+���Г��R���2�t��Յ�4�0c�:�ڲq�p:U S2�t-�L�Ľdm��J��o�,���Nn���T�*9�����P��H��/ɍ)	A���
<0�N�m3����$�k&CR���{~=D0d�?	��׹�nD���8x�wk�;���#8��ͼ�a=�EK����M�
���*�Q�M��ǧ��!�����N!�� �$�����q�:T�V��l�do��%��.'�05o׽߀����w�:�J�l���IS�O�:O�c�:S0S:�Ȇc��s7��G�7�1���	`�Qp�S�r[�U,�B+�K��˅yOCCk��)ਡ�6cz!�+���P��$��H����B�6��^#�:]���a�e�H���R8!���+�0Ǩ�Jϣ���O���En�T�]�t��(��E�Q}K�� �[��z0>N����)6�M�<����1)(0�$(6ՙ�9+�ְ,����-m%�l��ǎ򍙔.�ηS�,�i��4k��[>�w7_3�M����Y^VUv�����ڻ�(SG�튨�xEFI�5����]
Ə�w�;�$��c�>> �,����1��5��偭u�I�O��5�v	��G�ti9����H�:l�X|���(��#>22�Y*�6[��-�7|A������� {�'._5'��˜�|Q!N��W������;�v��҇�=۾�tdE_�0Q��2�-��$Q�u�;^?���ˎ�t�+�3���%j�?����f��4�A��*��#\Ϧ��O�"Ǿw6cN����|�=�;�5�mD�~����=V���_fe���Vͩrַ��6�E����V����w��Ev�u!�X�Ao���[�e<�s�a��^���Q�U��9 %նekJ�{�Np��yU���/^�����5�����Az����'��8mum*�x5ѫw�M햒W*�����qX�r6�����ƫd6�E�r���ES�]��N���2���#)�eU��V�K����~���>iD/H�7bO7˩�3�d0�÷��*�[���˫:��q2�>ì������V���o�������g(E_��d��{�3*YS4�Z�2pp����~�3z6J�8捬�(��N���7�w�ص��$=�uq�Āy9v�����?�!�_Ƽ��gn?y�	�����	����X�Im��,�(of�*E,��eUt��s*4ވ�Y��!�v?���@�C_�V�^����&��H�kM�ŒM���dQI��5���~{^�H�v�T�Z��W�� ����S�i��4����C�e�l�?�������E�g�p�=��v�Tь?j�O��}�Y���9���혛�}�������46���g@\lݭ�*A7�$Eߜ�����lhQ�|�*Ƌi</+��\@�meՄ����0�'_�5��f�xw�xʔ�ix�+
�k}�'v��M�:���;��Q����!��^��2z#+�jP�}"�f�'�H��џ�����-��!�)���t~	@)3L-�F�u@!��87gN�
T��֫��aCϒ�H/�{*qQ#�FNB�#C��K�K�f`�m�'""�e@>�����\>��o�I}e���b�R��J/���O[���8�����A�2�ϟ(Z �l��2+{ȥ&*i.$[t%��f�Z�1,a�!��
��6��+tsA�k{�+�4.Ĥ�ATl���mHC�
(��c@�v�[��I�m�m�6OjͰ��c;@������k0�
q�t󅯫dd��������^��?����$�ɲ�������rV�Nĺ)Ֆla瘟�iCY?O07�&���	nV��%*ձ?���S�90�oyy��N��	$%%��WY)	
��.��҈��$�
NȒ��z�9L�����0� ���D4��<�4���he�o/����n�2ƚ�I��v��.YbR�?t	�M!˃�%s�]^�QE�������Ҍ���a1_��8X��o
bX`by7���|�랫����@��;f�@s$�,���B4)M2 ��u���� �w�w�?G@�i�`�퍈Z2�M�7=�HF�4�f+�����`�;.�0�E
�ū�X�{����nJš9x�%@����.*�sj	�>�*c�B&_L;.Jۉ&\,�.-}���̳��n흖�K�zE�~^]�a�"o�8����;t�}4���F#E�.--!tp��������=�B�#���k�s���<#͸�e�U���������r��?ߔB�X����yzrː�q3ѐ�t)rP�"���@��������F�17�w�)+���l�����G~����S�7t�/>��a||�yz�K�u�^ ����wf�'�,��sL+'��NыyyG��T�Y�h�ҨK�Zv�J������>}�8��G0r�ã�CF������o.䜈0���嵱�#/K��[��@ �1�g��L�Pe���zM̭*4n?����<�*�n��<���B����|C�PSSox���.���]_]�?����@���@}�bn%�%۴}08q�����cD|Ā2�H2���<�0FT�lf6��=�E%'��yqƭ�M�1jb�C!`�}J٪>�6I!sAť!��Q6��j}g Q��Z�S.bJ`�l�/���R���X�\�`����Dt+b(t�����K<_l;C� �G	f~X�|�/���$A����eq�`�w�#}�S��eټ�КA�B�j^�l���L�@��t��))y0�:�'3D��$���;�J˂�!� ��|��7��	�{
�N�碚�IDщL�y|<P�n�ʒ[߶C�Jյ"ئ8�XU��G(E5�Dq�г����P��[#8�k�뫖�A�)ç����{%�w-4���^Hl�[9;a�C8~�����s���n,��&S��$I�K�ym�B�Ř��b��<O4Xf�X)��Lɦ�;N�D��G>�~>]�"���7�����>��t{������;��J����nL|8���uo6��o	�j.���uY���3p��I��Xi-�x�Vh}�y�`t���M[��C�����Z���[��Jg��;(�~������������ϙA��^.�W�Ϣ�ȹe~$��ޅsw�vp�4c��M�d����tδ���ܦ�����]�_��>z��9�39F������"�w�爫r���{#�p,�`����Rk�p�n~��z�UF��Cc̛æ�rlTE��s����;��}O��q�&���+d��2.���A��]���{�vȚ�{}H>�j�-gM��Z=Z�/¸r�������MR�1�*�h�����͛1E��l��{�kuo�i���}P2%y�����1^L��������z|��Z��Gl�ӷ��E�u�Դ�Uj�HKJ}���w�H�1|P�Y�������!!I���ޖ�<��}�3�W����+&�u�}��M�B���6���:����>D@�������Sr�s��|��g~\������|Q�k�妲�ȡ�!th��}�)gJ�!��L�R��x��D1����8��9�(��;-N��P������lf6u��(�ײW�^��>�j�ѱ�?�)K�zm�����WOU<B73�vJ�"Y��E��}���~ǜ�B`�4��j(���7!A��=sX�F�l��w���r�x�rƺ��9������h͆���OG�������A�
#Ua������� ��*<��뚈ߧ��I��eǤ�i�b���@���6H��R�ơx�4|tz�������]���I��D{��_sM�@�J*:�2�M��Ӫ萛�K|s��mݼzyz_�\�P����W)*�y�$�Ҿ}w8�oS�y�������;���3��p�|���r�Z��Xí�P)�����1�AM��ۆbHH�az ��?�����C�|{���E�jxՂ!�pz5+x�^>Se���:��V���IJ���ܝm�l<%9��<F��Ď���4za�L@�W�%����T)�n�j�?3�=F�d2J����g��JQ3���O�&$=Wۯ� ��l��r�#5i���0���`>L��2���i�Zm6Ȟ���?����r;]c���ϽC)fA��/[5rP���f^u���A(�]V�3��$k�M���߱dY��˽�P>{��>A*�Ggg>Cpl3t�z��jz=�/--m1������pR����tNL�a���Mx�|��w�a}ua@��J���gt1V�Ou�sЧ�.p��,���6�-6 �w�+i�zq6Y����@�{���C������>v�z�/{/�^�����[~:^�pa��c!=_b����]��;f|&Y�K��(w�\t�OW���} ײ�A��l�U�w�T����QA��2T��.�K��%�}�2 �@%N�9���k�K:�ݾ#Msf��s���Fڌ'��ݹ����|�س!�?�w��(��	z;�x�����Y���06_��v�cb@B�N ~���Л�GUT�~���w[���!��S�1���=D!�H �MS(0xV��k�|���	˝�tq�b�j)�>�<j��j�P�`1�<�Dy��xX�{
�h��>�<��[%0!:RR�;7n���F;�ޅ���dq�	��j��mG� �������c/tD�˱�Q���r��M���q^�;��M(���`xؿ�|! 3���I�����(�!�c��I�,��`�F��������fT�_��3ǉ!1�|�x�e�w����'���,b�Y2=Y:�(C�Aq�I����(�྘'c����w����e/H�$��`��{B���Mg���Rj�>OXђ0����E�b��'��8K�T�;�{V��x���U����!0�(�7r��i��!���+'|={3�i�i�Q��V��1a.��ϱ��܁V��b�߄���ӥ�C��L�s�,5�>Z�v-�Ǩ6 %�b)��Ĝ���\�� ~\���h;��Œp�ÜG@��Ɂ�K׆t��M}�I��A3������,�-�c��+ |OD,��{������ϲ<�r+M,�r���&Y��87IH o�&�\@/dK����e4�)l�����:Hg}wz�p8����u:��)�u�-^a�۴p��p���=p�T��Q��?}�|�[��UDDC���4Qc%�1N�x	����>_�n}TI�#�|���kc�I	�ߛW��o�!���`g� :ޅ�]����>���N�+��hv�v+�U�0�����.��cJڭ��
�v���<��$nǜ/e�O!/f�t���� Q\�b2����AZ �̟��=Wz�&XP|p�#��^(�h�9��7���Xz���cT�'���(�^O	o�J������E�U>�o�y������T���y �<���y�
�i�2��T/s�X:T��g2�=~ۿ�* ���1���kإk;����7R�{�3�����z6m3J����L
���$Ws�1\fֳ��.�㶃v�t�O6t�XI��dEױ�?��a>�8��G`x]�W�j�_[	z�<(<��0����Ò"N
\��I_2��r�:r��H��S����X����32"��-�}������:t��e�I�V2-�o��*�m5�z�e0ض��_��A��<U��w��)�%���U�_�(�=��̪q�~{1/}9�eII�Xi�]~�	�[ۙ�0���М�ܳ�lũ�fa����+bn�0�%�g�e���[ߞ=9vz���ήM}!Ao���>����Tk[�1�}����B�a��g���K,�\)���f����	�A���I�D�zќȇ�SO���i�c&7�o5ӖhZ�Z�Q�>~��4O%����S$�&R�=/9��2��ߋ�E���gW�H���֔��Gg=��ҫ��[lT3p�ܥbP[��X��:��$d�r�Qo��e�|��c���/�Ҝ����;�p9z�H��}��`1J��vk�qG��>ߘ��1m]�G��sj�<p�N���u[�}��9��Uۼ��H��Z����s�8�����D��������uY�g�v�E)X�9x�/@�ů����7��\E\�ͻΉF{������%Y��sM��D�ѻ7��]�t�V�%N��z��a�l`3���il��!Mx7kV�La�����Y'���'�˧>��ξ���XK�6H8��|���������48c���!#e5�����hY���%d�&��r�'�a����`����|/�����j���|z��S�M�.�
�:�Ay�)*�O}K�}���4ϗ"��.pt��7O7�����tQ�CQ������:�Z�����/]�N���즀�h��`.�`�r��zΏMJ]�T
ڣSL���p�/����֩M�n��0�y|܆�n�{�-�!k^�?,��|}3o)u�`��[�q/zAp�E��|/����i�nx��HyϕU(�ƹX�2����crd��]��q���d����u�h�F��� ��I����X݉7BqTK�����ϨD���NC'��|<�6�7\[��YJ8#M|�������T��J6d$��L\�hO��ҹca��h\|f�{,�Z��[���F�ά�(��_;d�|�y�cu8�Q�n�W�/@Q���#�E�������'�gs�Զ��|$����Rh?�-��b�ai��"���*v��I$�Q��ڗK�o���FY��� �����Y��f�����]i�j��0�ಝ���m"E�I!����Z�i=�{K�bi��4�e�T���6�))�ONp1���H�?R�i���o�(7������C�wD`oH�@q�=Wk�О�|Ǎ�z�1����E�55���Ϲ�o�I�Gi=!F���}B*�E�����O��\�,:�
�M�7F��A�kuzv�|��qke�
��4;h���дS�
�mz׾{ ��P�s�����D��dB>u;�^Y,�'}�jRz����1bD�����+���B�l�.ί��[,1�@�@w"��w��P��=D������;u���oN�M�V�+P:]�	(�'����C��u�q�/i{�1���d��956�3�����"��t:_�L}�ؘ��b1h�
�F���^8E�HLJ�K��&��y��
�����?���Sx�!ђ��IU�~�����S��-�I��ۗ�G�7�ׄ�ƣ�x�?���I��4�ż!�К�z����)�!D�M�}u(Ȯ�C���B�xV}�����-]n?<p�Tq��=C��������B\��	�/@�`0eͷ�6����/]�Zg ��,{�B_��j�?��"������υa-Y�l��GDD��/Ҹ �8�a]��㠁#ѳ�������g`��h��W��Üs�.~ܙ:+H�]������j���M|5qm�k����uc3F��;,+����3س�4�!<7h2uV�՟bA�KIN[�,������ge5�m\���j�>�nz0:m�u�,�x��;<���՗{znw�|�mY���	'&�~:E@�`�|ɍ�"h8�U�(y��q����ׅ������+�4�	\]sMK}(��.e��%^�~�T[�nRII��X@��`��Ċ�QyY+xΓ1�{?�]�m]-�X��k��j�����M"_n?&)�`1�W�l�Z��Fns��/n2��.�#�bb�uB������~�5�T� �Ic�����qqqՏ������?;����̂Pr�pl�s�~�7!�TOU�UJx���S��D�kA���C�݅Jv�Se����k���[Ff(m��7A������D>D͍������1N`�չ�9}�����}e�^Gk?|�~sl>++��}9SR�����Q7��z������)���1VUQ�N��B�M���M1�]�67�L�*��1(�Sd��Ϫ����Hu|����=��c^�oۈ���+'ئ��+�Nw��GآCo��()̾�tO��� ��	Vݵ��&�o7{�c�߲Ɨ�N���臨�\�	>K�|0|v�R��>H��Q���2W9�_�:���8*�gyxL��K{����b(V�2�x�Hs=������p��q��Y_q��M���Wg�#^�w����"Wƪ�|׃�o����ܝQ�x�I���R� �XL�J�M�~����d����s�+qN��J�(S��sc��9�c����$���!�]׸��O����$���ם�s���?D<�m~�1-Z�ߝ�E���ĳ����D�,HՍʑ��Xt�i*�8)�d�H�^r¡`(�9��R�@�㘏c5�S\��VL�8�$~0)=n�;l4�wav�P���d�O�����Ko��%����w�{���#��'�ܦDz%�#��QǝG�*9i�/����9z���U��)wwOF�Q�ƃ6f=>-�yD����q����Pu����D%[�(	��J��*Tӆ$T���A%-Fh�eH��l��2Hƒ}���2�f~�ROO�{�����ǹw�y�s^�r�"�R�(��	i����N?�DO��Q��o�_���諅}�Wl�H:6��S.g�.�;o ��8^�`�	��I>�w9}�k�q���A���s�y�,S)�������7���m�k!�ե�/�[$>�}T=֜)�]"A�'d�X�'�=������b�'y {]���9,���h�X$�0���'cMA�R��ٓiE�7�(-����rS�R.5�Snm���̱㓫��B�N2�йW�����2-%��A��8�\��L<H��S�Z;V�)O!�2��G.������������o���؋�.r��e]�J*�̍�ش�bR`�87>*
z�K�;w�6Ğ]B���9�H�c��p��r[�M���,��Q��ev�晍�}�x#��;h����X}��X�!P�����8	�
 �,��,N	+R�iZ�8�Ο8�xT������fl2$����aï�����׍$����E
��TPM}I�c15!�9��F�^:'NT����#�z�:�0��lE���
�����i�|���h���K��(9��EK�&��L��q���w_s��}2�J�|u���GW�6���Ls
�r�-j�l�u����]��j�=>��G!�S�*��U��Q�_w;<!h.���Z�.����@����w���%d���M7s���6fۆ�93��[�QC�/��fa��>�I3���
AǪ���~�b�`�n*����1���5X�;��l�0�@���s�����/�4M+��9�����`��G�rǟ���� �B\Q�򁓜`��i�j�C4M�O������f����8P<���E" U8)�!>7�l�A&#��R607���P]G��;p`�^�BRIM�C�6�W��:�O���g��ks�w����v�kЩD큄i'a4ݎ|$���a��������@LK�O�AL+� T��^t�/�e������Qsu�r�y����4�B��C����Z�v=q1���χ݈������sk�a���UE���`���$�>���������(��pa�Ip�o��� *T��nw[�AD�ʠ�C�;ߔ[��d݅�������d�:��C�t����3��1��� �zi���&�Z�%gY>@�y�ѩ(�K
���v����%y~yA����pY��]�Su��~��!�`�iT��Az����9�	n@e�)Q�z�&���樦�~޹�jE֌_��N)Y���:_AX�Z��(�'9Д�-^��5�t��q�p�r9�1?n���1�L�ٞ��q�S�|G<�����[��ek���'�<�ʁj9ߒ�_#�g}I��,���ʺ;q����g��I:e��d ��=9B����Fl��/G���Ԋ���j������p�pz *�=@o^|ɎN�DVd	���|����Dm������Di�J�(s�@��Ld_Rz����Vk4s��x�+��~W	N��Tg�����|�l�@A�Ӏ��{�s���x��*Tr�Pu�1̋��/U;A��S���jo �����5~���x⧾�����\7q����x��O��Y�<�=`b�P�/�O./�0w����`t�{�d~Z��5�*#1�x]c�]� ��2M��~���G�{;���Dq?��(e/��}��������?*|3�GT�0�ew��Zi�������e���`�j7������O����`�a�7�)9pv��<Z��<���i9�S�i���҂x� �U�]��z�f� ?D�5<	���L���}�]�5!{�솇lL�����Og+��7$zj̣C1eK�����4�{�^��U�A�-��R�kK+�k���rϽ�����!TYXN0���h�`�-��4�s�-����?OLܙ�_7��z�����H���ӻ���9%����Ԓ]5ks��4�9%�n�d�����2�o�B:���6�Eݾ��$�+w�|�l}��8�aE��d��~�Z�8ܗe'��*�>,�V(%��"7�q�%�"!Y][��|�&��R5+�\U�S����k�4xZq➨ΰ�!d(��/�ȧËki��엞0�6����=@\����Q5r��y�������jn2챂�����'V���qչ��d"�����=�Q*�8����1VNX?y��Dǀ,�"B�*�Z��;1�}�j�ӧRJVu�j�d��6~���2i�Ļ��g��XFу=�#�k�W�4��x�׸�
h�d���[i��)5-!p������F�M�wE~�愾w�ُ
]��$,΢�4Ŕ:SA\��k���^�gD��p+Z����C>��g&jŁ�i^l���}�G�/B�����[Q�����B�+����!�5��F��&�����r���wza��f/��m����.������˧ߌ��@)�����]���G��\�Ou�j�����Ü5�?'����3��LL�b ]��X/�����3$���$,8�y��㻗|Ga����"�l���.��O�&��*[����V�#���XX��>�~ $�����q�����}j��y��o��N}�� �?����G���r���1sv��`����i������t-�=ĳz�u�F�b�+�K�b�guO	�S��v��0��&4�ީ&M8d�mj5�*2eUH�TM�Up��a;���.��6yζ��ri5PHט�Rw=OD���oE�~ڮ,߈�R��6�v�9�~��v5�Aj�<S�š*����ش[N�/���ܝd�ضT����������g���������$��B�Ŭח�m��*�����}�	a�b1�qv�M�n�uR\�e���.g@���R�U<G�y�5jv1	�M�S��|ب��E����S-��ȳڴ�=.(U�7�>��B���b�($���m_������?q�3'G� �
z��&��Ld��U:�6YH��Xv��(1l�Pg�CߥW�G��2o6�k�;�8g�l�'E�S�s���DQə�>���g���o�T3�H3�����6�H���"�OM�q���O����N�������?*!�t���5i���=;���`����r���kb�	�*�H܀�����c���W������7��Zy&J�������r� 8�OBT���8��D���N�f4�ӊ(��=�6���K}��~��S�����:N��d��_�Ui�{�sb;���1��B�y���Hpb���? -�ʏ�%���&`�'NM��]�0رg��E�i��b^Ӄ8�;� ���g(����4^�zP�	�z���a�i>��+��j��L���d�wt:A�?Jok���R�B���wg�H; �5خBf�
��=F!�Fv�"\Z\��߽.�b��2�-��_&|�2!�O�����Y����F<�9I�{u���8�@�"VC�J1[�ˇz/3صvQHW��l�4H��ރX�ܺ1[�ɘ1��m޲��Io���#P.Z��9f�0�lSIĚ��]��F|O�G�I)0���z#��p!��$����'��#��<��-���T���K�`������xY����<�6�8�yzq~�7�
���jf��W�B�C!R������S�B[��2�3�����s���i�5��朴�Y>�C_KC�_1��:�'f8QHbSM�5�]��O
JrΨهѴ�����A{&�\0��#��V�; e%k5p���lZ�PQ�ǘ�����FH���v�������R��O�Wq�Җ����FO-dÑ޳4���/�L��i���m)'D*��\�����(%D�_���gsc���垀^�zjP�����=��yٴ&U��!ϫj�4֧��[:�Hm�vE�q�=��y'��$�����	�%y(��t�7%���c�����fϘ��>Ru�|O���7!;���.Pə��Q���1����fOL>C��øI�� b����LE۩��x�0n'9���Ge���
eG�-�z����G7��=���)I���{�9�QQ���+O۽�*mW�V+Pd�s	@�vՈO|!�'�������ׁ.��w��<]��p�$�N��ܯ�
�쿣�D��_�KU�R��e1����{��Э����w{�����m't�����E�Br0�}��8�=մbnO|�@���Y<���W/�q��~��}������w�+����m!h��?3g���
��({~F�!��G[���ϻ1�J ��h��o|�s��&!�#�
��9Z�ýd)z+��P��,�������K>
�`[ˎ9���/-/����áp��P�[�����7���QV�k�<��(V5W��S�[�IF�(�$f�C����>%�U�җ�H���"��.	9��2ߥb���Rz�m���x��oZM��%!0c�.��|����4��ͤ���N�����T�j��z`�.��	��s��ɏ�K��z��7��gb>-ut:����#Y��5����-�_o1A�R��m����J��1�0���������_��_�y�|����{���Ժ���d_$����҇�t{RW�S�+i4g�*�����xK�B�!�X�%� � k�,�(�Q4z���N�iw�-H@��J�4-�ٓ���A��w�8���[S�>&�:����o�G ��L�CW��v��d�7��A�v�Z��]�:M
,t��U��w�P����K���6ᮐܭ;D�b0co���/)���$ˮ������I��#�j}_��shE���A��L��}�9E�ld�S���i]#sȔ����^�8"��v4����,�����#F���%�]zo�﮿��A1�U׃c-�����ۚk�yn;2'��QanT~�+�r��������J�6�N�V�I	Cx8�J����q)u�x�cH�6ѩh>�z��Fȭ��1��#�e"s&��'c����c'��w�4uVt�'Z΁��3�N,�i�Iq0኿��-,Y�x�+s�*๪�HN7���2�c��%{:j|?�O�XKwh�������q�䜇�H���D��#9��ƭ��<ӯ%և�6%&~���@2֪�f��*�|+�;�
1{&��B,�* �f уf�i�~�Y$ }��p۴�h����@�gW+n��*���ёx8�>kB��<Ō�i5��ަ���O̝���\�c����2t|��5�7� pp�^���
�h�tp�m�H��.���%С^�S4��$���{������x�C_K)�����.�}>�u@���f<�B<�g�*����%��u��ؾd��u#v̂�87� 4$�z-������Q3~�ѿu�NF�.�Y���*k�	��*�n5��GQH5�T�b���q�}"v���%O0�~M^�[Z�qi���_�5;͑���]J���'���L���8�bcp7��sH1��4���צ�@��`["c��^����V�M�-և9f�PTQ4��@�T�LZ���~m=�i���Fy��7}�j�F��A'W�����W����'���H��xN[�*a���%\kl���;�r'"H�UgT����<�	�/�3�F�$VC��c;���
�����W4.��2�!&8�^b�<ϜǱ�GS{�㨙d͇��_�JAfmF�)KE���d�e��o��=��$"]��ӹư!�\+$�	abjnw��2H��jU��Q�Ew{���v��K�r�����=+]��q2�ys�9��1O68�uz&VCF]����禡�e5�him�W[K2ϦM������|�_� �dp�N�Kz�OX�����,��Ko�S}������S�VG��^���7�/܇a��v=���SG�> �(ݙ�`�:1�cv��KʰՅ�n��Bj���3>�������_�7ls���MשM�h����e;�q�C�2�g�>va���}Y�gv��%���2EEk���8�j�����u�EV��tFg�[u���A��y���Sqz\E`�+�j^�"x��eK}�j������������'њ� Y6����w2򊽕��ȳ���J?>�����HN��)o�Ɨ�cmF�f�V���(�;ĉ��d�A8�n���hŰ���]��	�ɇ��S9G&]d�^�"��*���H�+PM1�A���)̀y7�y%�ܝQ(hu|�����F*�F�����DG� ����V1�����y�*��>��^i;d^�y���S��1<���>t�_i�#h;&��CY�ċ�~'�����gT�{�RW�m�]St�?��mxQA+�J�=!G#�u��90��ρ��f+��y�vsBL��Ԙ��i�G��=��j*����?ω���%(\:x�(������-�M�=]u���$�R&�Z�]�]��c!�K�����שD���u��D�U����***����1�݊�-�/�ݨ��� ��
�./���&�y�8A�L��|�L�u{�Ǝ�����q?g���;G��>wEF`�pq�+.|�?�n1v�����\t�Ͳ�*�4������LHH��(��읬,O:X�G ����ÿ�����3��Z9�$�/Xm������~���muQQ��rD��Iӯ}n�z�S�����X4�At�������=8dؒb?S�����Qd��p��в Nmub�qή��E���$�3<�36f�����N�GH��0�^�����;ٮ��AX�w�ݯ�q�N���9�}N��d״�69�D4�gL���H=%�N����C�8�L q$}���5����������\'M����]>�v�"�x?��G׿�+�y��k�=��V�[�h����>�t-������Ih�6�"<Q�\���F:�d�0=pk0 �2���t
g�!u�۝����1��=p@tqv4��Ǐ_�e�|�H_��,��)��������)������X;X6� �WX�S֜�((�p�����
�]ݾ�O!!
����d�V�#L��"a<jFOT%~�4.,£���,r���ԫו�\�b���Xyഃ����E�¯>gס�ۦbjιf�4%�ڳ��|��\iP-�FjV�n��ɉ����{��I4 ��u�/}���aCO4 E�]?{l�H� ��Rrg8����OH�)F�2� ����j�l����h�]#�w��ߺ�RV�[.|� D&�tm�̱��خG/7��?	\@���p[��Qz�ñ�pZ�(�"H�&���/�5腌z�m��_�v;�
�"m����AP*s�9�Fs��~%�⃴��D~��;��h��h9���t���7O�	[Ӆ�]{�r�h0�Ƚ� .�ҧ�'���ÿ�k )�����f:�����'�ک��ls��Cv9mVh�K�g8���4Ŏ���N�޼_�0gl �_-.'�k-֏�^m=_�DUљ�r{!���=��D�y������-IA�V5�V��(���ͺB�]ˠ��m�AHt��o��|�*�B�o�q�)Fs�S���\�a��#����U��^dC�}|�;xT"��7diL0��l�[V_6��_�F5�<0+9�<ߋa�XfC�{��<A���*�:��zߎx$3G�߰� %z����61�m���H��#4�k��Zf����� 0|�?�L��z����	v��z��=� >Z��,Oy����f�h�P�~��ך�GT��L����_r���g�3�ٳ��ɄF�#U�0w�4\	�sk%�b^��j��9���bC�"�����&����c�����C�-v��b?��#o�T���\�}ctKj]�������7��楜�0ȍ�Zn׊_'%ٖ;:.s]ab�?1��^���==7~'����`\*<<�x��.?d�p~�O�9��%�^,��|���t���\}D�x�[�17A<֑�@���l�����+���������փؤD���)T�&m����!j�yهL�<m������Xu]]�(�� U����w"}����mE��KX!�;؜�'�w#f:l�t&Cc�����CO͞�&ܐ�����Z�����F9Cp�u�s���+YN؍�"e���~�m�bZ+yk�ß�$8�Ϻ�O,M��@�(%�	zY(u5�V����Kh�茑]��'���U�.9Fn�i���?���Ȃ˿� '� {���~�0��X��͝�ps��c)�T�ݻ�w�F�����_�a�C' ���H�������� ���$
������iE7A��+�Bn~,��<�{w���7��M�]�8��ʦT��n�����b�밯!�԰�H�-��@;�n��AZ����1d�z�bI'2d�&�ow�h��_�#�o޽ӭ�D�,3N����S�3���s�0���:��O�ߊuƎ��ؑ�AP�������e ���J]I�
$�p�V$%Ih�C�# �l ��0��4���ς G�4ð�S����k=�J"�����9X��Ma�$�m�����`S]�r� �ڱ�#="�Vy'�������C�&��#�N5]*���|n�>������pVf4{�N�m����VT�ȃ�@�j�Weon��B�!�W3g6V��c�������8��*�w���D5�W��g��HM��;5�!2�W���"�^v��'��<�ʎ�}���@�i��i�jm�y�f�y�җ+����b�Zp�pN{��������w��o��yr�������@����tO���6���xŢ��c�fj�
��ڿɗ90`��"5���ަ۲��5��Pg�Ma� �g��懷���ܛg�Rp�־�<�h�m��SP�9��~{܄��#����	Eב��y����>G�»�a�FFn��uZ2>MA��,�D�.,,�?��jG�aL�pK�)���9J/��c[&}�k1��D����Q�l���"�ůI��Ѿ{���K��(����3㝆-�f�9)�,�3�,|~0k|�^xxx���H��<h�#lO�s�F��FA�S��@<�|��OZIIi'�lB�a�`0�b��Ν�FT��H��;O��8 ���c�Y6Mc�Xy
IÍ`p�8����"���� i27F�����|�'���Vv$t#$��k/�k��:S!�6����	%�{�+-))�R��j��|	�ן����Z��_lYfl�h}��>2�BF+(�ӷnݲ.+x�pp�lҰ����U�?�𵃠�H�BI���6b�NE(/��F� �����?֏�ؽ[��˗�&�E��T��<�}�*�c����2�����I"h���&d�l�Dg�U�y����Q�b��D����]�����M��f�㳁M�'�D�\G�ڔ��Be��X��:{��m�Ȃ� ��
p3�z/e\F�S�}ς�?>�.-#&N2�0%���~H��o��?f��e�'i��.P�	����l�rҬ��x/��D|����jۧ������[�K���o������n��Aѕ��+�`6�T��xk�.�/Nˤ��b�>Hj>��Ъ�Q��t0}ͺ�+�p���NF�`;���6ӄ�TC}o�j�mM{�S��خ#��	�d�[lRg�+�[��r��
)��_c&$Jͽ._�A�*�����lBg�}���O,�W���o�8�k��ȳg|i~F�&$�Kb.��s/����B���\�������4��J�/F:�����G�`c|��[�YC��˴`��Z��鍺@;��ȳV4�UOZ�w
�X�΍/��~��k�E�<Ԫ3�\�Y���~0�w%��a�[W�Au�VqK3�>w�M��t:}�q\ ۿU<�ƹ Ε�h��t�L���n��P�g�p��_�s��j �y���c!c_i��r��T������<R���������������@N��`*ԸĮU�MW� ���%�w28�Q��1hb/�; 5Oo˳��zC1G���'�	z��4�[lWc1�u�U1�����R߿�8�-�4�0ʺ�i�Ԛ�`�{�+��b��̿���{��TTA�Q����\�G+<����8"j���ʯ`�� ���9�����p}�^�&0���\|!/jtM��ᱬ�=�-xF�G>�����E%� �+��W�P�@8 �X�TJ������r��>k��5�m� �[�1�� �O ���̷���Y+��b���7��>����NnX�v��i˶�������-�,d�'��YwQ��R�e��)�N3������w ����b|U��- s���?o\:�����V��'s��r��e�u9�zd=�p��fiM�B��/�֢u8%���y�pU���_5��_��� 	}8���6�֙O"�6��{$ X@¡���Q���m�H��y�̃J$Cg3�	�o	^�A�������ÛWK��(T��G���D���Ir��� P���D�;���	`d;�+z�,���G��Yr'S!�?��Z�U��P[	�|��E� Ci��g�)8��ދ����D�/'�����p�HR�0�mJJ��ӧ�V��K�I�vx�������~ҾD󼾾Tss��P�K2��2�?X�~�˦�99�ƹ�#ԫ��{�ua�.�;�j�e�Х4j��D�hxW�GUb����ƞ�ȼ����{S�Q67�c�#��e��+�^�S_4����v�����(�0|r=gw��%��1�T"r��/3�-j�'cjVR�Q���A=n��i��Օ+e���E-��YlS���֔z�}���t��	_ٰ��<�l�<U��&����z$f�ovpՔ�����e�DoI	HG�2�x'D�-`�eZӨ8&u:���vNx}��F�����Y���P�
BX<)XG�9��}�.JER�����<5|mh�.O��aT~�,H�/��x��*���gv5��T7%Y�̼5��$Y!��)���'o�׹�gl�(a�Ay��vBŖ���h��^I:5]l���%}�>�x�̓�G��T�6 ���I�-�n����w��-�.��|葽�r��j��ؼ9�`iY���ܱ�����[�P؄5�G �d�7)�t��܁�xHT��Ҥ�s5��ψ_����(ڠ��"���=��Ի��l�܅���޷�J&��0��G<�����p��;��G�t���>�i�jZ�nRÞw"�߼u�`8�~��k2� q'�~r��Y�2g��z ��f��/�?zb�{{�2����ڹs�ѧ�P<��>p������AW!���R�P�U�w!�w�zCH�����Qh�	���Y�z�>�Q�E]qk�tj�7�n_F2/	�Ϋh\�M��k����+��J������"�-^����+�s����0C��kߝ��0]F���d�n�����䪯A��������O��Ӵ������~����{����z���P���i�5]�}KVD_��tv�D��yeT�sF|]������\��L'�j��ɠ E5|H��n��ڐ@u�P�����70I*��oE���a߭�@���&VA���FR�x�9�U��[�L��m�I����H���C�9���{V[���Qk�"9[�����j�;99��P���$�����=�ƚ-ym�fZ�i�wX)�knL�u��ҝS���2K6&��3ɨ���A9�x�8Y!3�G�#����d�c��m��@�y��{=�)�y�������-O*m�l��z����Q��l|9�Ҙ��ŷa�H�$Q]VR�ō��t9Y3zϻf&)?�Qd*�����䓣p�\�Lm3��
�x1.\�<R�]U�5_�wU�Wfx���
A Q�	4]a�^��Dkjp�/3�p_����WM��D���pj"Z��������W!�8��q)
5" B��R�}�U���k��Uy骿�����r�6�]�I�j�*w����y�W�}Ej���Ua�R>���ٳ��h�Zڧ���:��ؑ�xy�n��vY9���3��`�׎��/�7ФVK͋���XD��_�A��5ر_B����]�/�̪`�0am��3k#٘�5��B����L@��D
�\�:���{��7i/΍�**%��"�kTBqG�v���Q��;$�@�o�v���E��&1SJ����t���t ��Jkg��ר��0��Dxu�L���������/%��C<�x`�G�?}�6K'�3�����FtN�ŷ����oWpƔ{k>�M-���S&����a��և�]y^r�Gw�2��K?o��I!�a�"����Z�,~z��?����D���>�ƽ��]���D�i���I�����+X�Z�P�Ļ��vC�H�j�z����mE��eI<�s���K8�:��m��1�y��>�+6��zT`Jzw���s���[*��|H�*��&��U��q��Jv��V����������C�1�g�t4���m
�`���'�O�<�_J�qs�̱�΢�S�2-*=�|{~g�����z�b�x�~航x^/�<����i4kl�Γ�(�Z9�T�-�Y/wy�a�­5�PP�$��N\C�b�s��_��8x:�x՛�x�4	��$��ӧ]'�Ʃ�M�s/�ٿsxjx���|0�r�.��y��¾7@%��eό�~I�M��4���x�m1�8(��<�{�=�?,+/Ox��ի��7�����8\"��2��g�l�i��"�ӊ���lש��%lD�7�Zn�68�,@��2��k�hFB��Zs���'y��~���w��7 d�>_А��}r4�OV�(�'�d�~R���d}�9~��V���c���|֞�|ㇹ{�r�Q�k���*�}#��N���h~ﹱs�`8etR3��n�J	|�h+l�/:3B�[	4��~T�V�W3��C��N&��"�b�y���{ϔ+ѣ&���6Xt��G��p��yw�QW�j�΃���kK��~�{bZu,���K��7nF������W8�*�9o��}?J��M����ܜ㫤��aVH�$Oc3Ü��I�dN�DK9f>���`���Ӭ��.�qC��h���y>�_&�1�,��B~�������M�9Ѯ�)I�WUA������؈��/_����Hz��H�Ϟlt�0l��XO3���)����ݽH�5��b��zgH�\�m@cǷ�Rf^A����o ��1�
 �$�a�/��"@�n���J1v�me۞*ڌ\��ώD�!� �I��W㊏F_ysHx�+g3�Wԡ.\��b�7�a[�*���D!͊�O��J��F_'aZ�h5,��ئ��o�<�:��'��٘"�T#u�+�w���=�;<:����3CTTT�>��t� �6A���
u����U]tJVF��?��J�2L�J����x3^���zo�C<���0�|�,���룴$w�']�A{l�������D�x4]�RI����A��o<�j�g��X^|������4��	�S␶߯63ޙ�GJ؂;�CAD������7���� Χ=�#�T�������g�o��Di��C�Y	En|۔��fZ�W�ߪ�pi�@��߇����vSsFfo8d2�5e���]���Z�J�c�#1��4�.�:��X��-j6v���XD�Us�3��޸HPX����PAŠx�^��d��*9�C�۸�iӦcQ���v�9^���g�ĝ76�n�Ti�wMv%3޾y�ldd�>5Ӷu/��$\Ck��m�#����(ߋ�
��ʓ�MA�b�����4��[<+�7HP�L-+�`?y�l���kܹ߯қj��}�wE�B�U�^��������G�V��w�����v�(��o`�x7��=ښ�Ig՝)º}$���	�kBEޝXep��'e�#���O��'d#bCC7�N�F��S2����\bl����?G����x�v,!�9�Z��TRO����\���{����+p��۩{=���F�p�;�����2��=4��r�q���ƺ�p�uI�SS�^��KX�/�@n¡]�M�>g\�?�69ٖ���l-e�0MK�����oE6�U�z�}��"��:��X�ij�E��
]��W��gO�uF���v�_,ܙ�8�5�-E��4��y0ͧ�zp��u&�m���u8�N��-��:9����nj�dk}�Q˳�����*0}{�1}��v6y�$T6m�a�OP	����B֩a;�����d�'��?�dpo�[A�4"��"������#<=?/>��R8}��)�bp�#:܌��'-��-���a�Q��F��8Æx���Tأ�gJ fQV�������'z�H|q�6�r��/K�Es/�hч���r�]G����!vH�J�9?�Ǒ'���}�{����\��iR?w!d�����Ya%��k��<ء�l�>o�e}j�*E���{~"θP�d����7iyob+ޑ�p��ҙ��u�s#r<��1�X�o\�FK���L�'�n�.y�-ƏK���({޼��Q�]�>�2l���"��;g���׼�8J/������k�
�&ù!껔g��Ϋ�ۛU1�D[��Wm)!F�H��J�>�,�z�����P1���g��8։���R�nC�*�](��F��:RĘϠ����/v&��m��t�P8[�	Wt�y^�D��EFn��Up�B��ʙ�j����CN�h� D�e7;���`�l�����>'9�\Q�BعS�R��Ұ��������m�e�^�^kU�{�E�t��In��7�R�^7H-�X�Z�����o��j�77-\B RخM�o��7u�=-�|�]�F�q���{�x�2��oߪu��G���,Uΰ���[͖�Nq9�ne^�3���$����n�"{��&{ଌ�pBD�6)np����P�}u�f�%6�Uۅ���+&�7�;pƝI��e��t�>�G n0���mR ������=��ه�^D��33-fk��>M,#�ٱ]�z��
�^
B˹:�O�+e4����|0���VnW�D�C��:ŝk��gl��N��Q07��Y~�YPӥ�
x-���.�D�>O5�W�,��}�L���Gq�O�C��N@���?�WC��Gvp�%G����M�߹o�qi���w���9�)*{���<����w�M��0��ќ�=�7��`E�{o3ڤ�=J	u���M����`8�By��~�r�@��Io��FeF�	�#c%I����^|���]�Zƕi_��zg�p�k�7c�{�N��M�4C���:Hp�Jl�˕�� 5��Ƴ�*��c%�|Vq;�j[��'}V��׻1ʨ��|yP��VZ�⻙]r-��]�2��M.�}v)�M�p��e��}WΐL��k��8)����P�"zGs�����T��{��e�~D���'vP��ղ��8�4Ȍ�z���U���5�c�۵g��W�B�c�*��%���_�N���x4��T
6��M��5�������=� ^BT	��S�Ps-B������NI��hD��J>Z27W{o�̲�����Wo�Z4��Ƴ��=:���ʍ#�C�J�"����hM����d��7$XÙǐ�}��aV�F���X��,n�&ڠ���@}p҅ �tQgS��`��/f�|q���{l�oNB�oB�Wr�~�nc�gE�RQWW�'J�q2��Ċu�{�|��|��Ys~�5G`�#ќ(�h#֟̕���{C|�|h�י�<>t5~I$3����2B$�C�A������7O��Qں�@�;���Z��N���vy|�kE;�1���2�Fq^�Ҋ�]�b
�{�q���/q/v�襅R�L̏E�v�E]�땛�+�h~��D�˟)9��՞ɽ���4��bU�Ç��{E@П�3���6��f��#�E��#������i�1��c�DR�G��%�}���>���.��\Vٛ�4�dR #���[^��?SG{U�-���0���YL�л�\;Ğ�%�^>��4Z��Dm���%%��ط^O�
�{��c�� P����G���ia qI����Y͇k�oT�l�`��@6����;z/�����]�8����6��G��l��TW �Z�Td��C�[WJ/�`�e�?�'n��#q���U�lÿNə��ƘaI%����.�}N�Jŀf�0�,�j���8j����E5�\�
�'�yf`{���4��MG�_@"�~+���Lyvx�|�]��_p�0��l����^���3M[�i
����P�S8��������j����{KCi�BdM[-�MRl=��@��|.R�r�U�����b��'9}f`d�}b%�\%�Ѻ�'�]�U�����O��:�����2�ڣ	~�F9IE%%�G��ß��'��Խ��|9�=^��+�z����-�
B�U�`�}��|�r`Ɏ���P?������W��]	�6�醈���+ƨ8�$�y��I�j��h�8��N�5�d<?qٍ��۷�:ٸ��3^%�BU����"!��|�d�vJQ�f��O��+��B���uH��8�s��s��`*�(����ʾ+���v�~�~=�ߜR8o2|�̾ؒ��w���x����>2�@�<q�Jn��p���2���B����x"�O��
��8�<N��9��]�T0�mlj0c͚d|�kN%Lx��w�Y�]��E�J�Cj�Z���7!v��� �d��z����5�	ԯ~�i�������y�9t��y���k��]~Er��YK1�e,3w�Y�T066ݥ�f$����O,��hZ)���67�T�������Z-*�v�ᾳ��$�{.g�|&g,�Дx:�����7o��(�WV}��!��ɨ�d"4�.>_�i'��,�]&b�n ��?�7�Yd���Z����e���p޴'�$¨��i�ǔn{�<n��%`i��=7h���w���B�ٝf��7ҩ~��
��aJ!dz�ۚ-��m��֛��X��KXJʞ�ܕ�p����#�QW�d9���
.��#5���j�ټ:2G֑�wD:T��^֗2��Y݄^w/W��-I�	�j�H
�BsHѺq� ��]�5-�m(��))�m���f�����
�"_r��]��N9�8���sPZ�q__Z�vZ���Q�r�0�kNt|u���b)|E��>$�9���s%QMg>^�'��=�-��S��I=�08�>m���
�pB�c�"���nZ6��F.|U��IJCϗ��-V쟝��ibF�D�#pxN���c��$H<�a�5_N�ǵ��G��7���=V��#^׹Q����[��+7���u�Ժaf����#VP�d_Z <a�Gj{��q�������'��I��V�/������ C+A��Ḯ�q�K�Q{���32|3dٽ[#��^
3�°�w���������wB���₵3�G��.uu�mI�{T��99¸V.U�Ec���$.mIY��l��Cż[5k[{�P��a�c�acrV[y�9���JT���>��777?7	�$[��䕕+�}���� i�{.uHs>[EE(�o-�6���\lF\�	��T�i����V��m�NDpf�����S���)����0
_�h�5,�8�4$�ZҞn3'T�a4E�Q�� ~�4�ǟϯliF��I|K ���2l�n��r�,Yŷ"pS�g[��^q�ɟ�"V�f''X�]���@{���e�|��l��Yڎ}�]��?��;��l��#MT@:�  "]�DE�� �*RC��JU�Ԡ���A@z�-�NBM ��Fg�Ͻ��y|I��k�_Y{�Ms��%�to&p�  �Q�?U�K�ו���-�0��$n�w,|�Gި^z_�O�֌g3�c���lc7$(��������6,�$��������j�
n���4��M����,|�ڞ��:u�t�~�!Y��A�"P�P�C�!
 �GZZ�h�o���f�x\g5Ϩk�8���L��}�ܕ������ɓ��
��;zz�޾��(z�!�_�u������!hP���>[Wc
�.dhxͺ-�
b�=�l��Ө=h�w���+}}�=�LF�5�X�xb`{}���xl����f7��P��йR�����3����>���z������p1X8%�5�O�i��g��sM���$��~�j���=|}�Ey��Q3ް��t}1|·)�N��n�<\�If�|ôN���:Bx�,�+Ϩ�
?g9q�W�\��z���+û���M��t J�NP��&�n3a~�7�A;���s�^G}���I�n{Fo�������-���<
���{�������6���\L��x�Pj9]����O\�z�p]o�#���v4��E|���>�]�7�ɨ?1K�e��0�*�8�CȦ�V!_Om�����_��Ѵ�Ut\i����>c)��|�g�G���W�����>9��*�U�GE��5�i�3:�xT
8r�q�+.�kv $��h�\��"�aw��X�x%"�1G>!�]ؓ>y�s�܏>���M���8'�)���T9���UZ��Ô*/��w_�n��%�tI³pu,��s����|�tީ�5 �0�ӡlM�s�F1��fߞ�� ۻO�J�����7�#rS�cSw_�!����N'fsE}�0�N�n�Z��P;!)��8�:�FN�הxٽ<�-!t��]gnW��!i�I��}>�����}��$��d����ʒ�`J5$%[P,���I�[�v�����}����޳\�,�.�0�z��\剿1����C�����O1���-��5;�Fn%¦Uч�S	z��qfPܡ"��3���F�y9�G&am$���mV�|�m��6r]�l�����\�b��!�9�������̇wO�N*�9_\%���*d}�K�����$2C%*>��iΨԶ����(٭������6f�C��s�b�G��1���4��<���
WO����~΁l'�t�N�F�-~K�G�޲:�KA%�����RL��u]� �,sݢ��*t���F�jPd��v)	'� ��s����T?>gf���R_
y��P���cU�,r��L�Y]60C\|�,ę��N;�����O��4�c�}$�H�+x��h@�Z,�k�l���U�bY?��7s���S3	|�^	���ɴ+�K<�^MG����-�t)gA�����s�R�ܘj�H�R#~ɒ?��@�s�ï�CZ���i���t����)#COiUh�F���p����@qK^�;���:#��M��D�G�oO8&?�µ˔-���O��P	��}��;�c�I�c���BUCF�A����W��dQr��\��z"dR�'ľ�&��!������D�y�yj��(i+Z���@P�C�Ů3ߴ��UԊ���=��/+���G����CyG���[O_��ы��qzV! ��):d���yH��R~�2�ϴyC��&
g��C�w����x���q躠�`^BAR�潒�;��%�P(g��`C	"4):8�G!?K���cc8'�?�=7��~��^��(/���>�=I`|��<�T_���`�^o׏���
�WI�Y6$]��F����a.)&Vj�C�ڙF5�c7]��<�c��T���u�:?�K�O}Iװ3�UWǟbѻ_
�!�g�;�t.���d1K����ɒ� �� ������n3����6ښ��xlu�\�B��!P�?�AD�D������n�>嗠�r�\��������WH�G�NI���
�'V�i�I��F��t���לP��i��_>J���g��'˓�OP�������+�=V7�e7�����e���@��-'�}d��= �V
`��Q�;T���)��˷��f`�y�����V�7�D<i�h�qyRE�Ud�~��'69*P�{/�Y���!I��vuc�G�M/2+�<|��-Hm#�	!�����������Y��\�����3�(���ߊ���.C��c	�i�e�J�v��C��#M?嘾�� �<��z�i�3�Se��u �z�Ǽ�3�H>�>��̯��[B����%o��x1�/�gH�Ѩ�h��(���Z�'�\[XLE�6���]���_��]�BI�s���b ��@~�C�o�S��X;���&�܁�����Ll
+�σI��f. �j~��k��ҝ��	d��>ᢑĘ��7]i� �OO1���ȼ���s�f'ţ�49�x;��j�5�P��!		�c��e<Id���4�
����>ؙ�Y�m���L��mO���#�E�)�(M��v2�^� bb�`H��'��kB�-�6Zu#��ۭ[�F}!�oٌ�vyii���/��zGs�f��@���	�@���l������C��V�����#���ӥf5^���nW����b+��&���e�ݗ&��z�t��gNw۹��}��o�rk�I�Z�;��#CEɯ�nl�'�kk�8݃�]t��wU��w܋�&coI䢽���1��V�9Ze�M��=�5��z�z��I@WUJ�H&��0��'�X���ӣ)��� �Q������k�qs����&ȶO+��B �J�򽀸������ ��������o�~�,��u��(=�4���h�)���M�U����d���IF]����Ȁ�4 ����'�LY�]}|rk����d�!�A+l���3ͺ�[���|�r�D��ʹ��r�X��۞�?�� 5�p�ҷ �0H�ډ~�D�r��������fy'��W9Ϡ0mANs��Wn;�A}��������I4r�}[�1��5�eL�0�`o������wR�gR4�tp�r�<�Y�� �{>�=�4K�㖐�E�$q��.�䵽pL��DZcB}^2��r�_t^�6��
��"C���D<
�� �|-���a��Q�M�� �n�H@&��[{�d��?�@�<�|��p����y@�j��<�^=DмU.���������(��m+9��K^R��H'�s$J�Q��/�� �B�Ul
 es�xO�_�Rw5�d�p��B�	��_�J�F�Ʉ�q�fA���jNv� �B�.K��w�<�Ϩ��U5G<>����+��m����" wM�i>& �e�=��ᇛ��u�9��,��J�7�A��eܧ bey�O���ݗ.�6s77��*�ջ��3q%)+�}�aw7�z}�"��9�Ol�7��C�<b����t*��@��ނӟ��M�ޤ�O�,Fl�a���O�ܣ^�R�.n���6��3��X�UH�*L�j������*FN�P����`f�9w�_����l�2t�E�$�f9J35R_1]uSx�#���8Ey܁�L1ں�|�k�a�n+�7%�
���F��'��,�K���P��<֑��-@ȱݔu��<^�tQ��w�Qn���1���VxԈ���"�&�G��\H}�E:4)�IDWu�����vw��_c?��$݉Ɵ*��V ���x��#�C�l��u���������on`t�y��D��;���cP�1�Nc#X��-��j��x�����S wd�ɾ/3;�|#��(���j E�&�0���K�02k]��4�¢��)���%�2ȶ�YȔkMD�mO��nE֭�r����w���p�$��I� e����[�R�_�*x��'��l�Z����:�#�5�9��������q? �6[뛴�$wg�u	��AK��<YLx��g(;`�WҸ!���Q�Y�0.������D��rzy��T��\7=Ww-�A�K?V�0ۏV��<Z��L����9:^������d�[��ք�
�j8�+h@͂'&J�⬳5a��0�+���+�d�7����I���a�,��V��T�}�nb(W:���_�|ч����ro�����1g�I��$5�௃������6�Cc'��iTF�iPk)��>9��pޚL�b�-@?'�L5��9�iHGſ�0(�;��b\��'���=r�< �G���� ����S�|t������)�ٸf�Έ�G��2�PU��������儤U@�X�C^}9MXmq��h��w������Z�V�OHх�h����������P�1��k=�@P Hc[�I�m;I�]�~?�z��N�4�N�uQ8��/��.�\�o/
}MQ�2聁,<p|0�{��a̔�Or6��p�/���&�T���~̋^b�Ho��ħ�Ƿ2��T'�4� �FI�+�b�F��_���ѻ��3��\R���>E���'�yn����^4j�ɲ��k���*���e�5���H6r;U���Й�=����� ��%+���.��R�|!~��+u���^~���q |��5�	؟To�n�O�+����@�݀Fɬf�a{YZ`V���G���7E��"6:�� Գ���n�"�om���	$H��ɛ6�
�S�>m!"auT`��������=Y���y2�U��Ǵ��e6��ڵFk}=z��@�[S��*�p	��t�%�o*�7Q�[N9�x�h�,0L�����d�W��E��|�r�Ԟ�.p��p�obz��p�@�o�&@ZA�Ǫ]b9�ʀ"� ��M�ɺ�}(784�c��!^�j�J��kg��Z��Ϲ��)���j���@�A�9�/<�7<6�g��燨C-���Wɚ�J��p)�$��񝂅���$	�q3�`'�ܔ=�W�?
y��Q���Γ�.a�s��0&N9��w^]Y���4� ����h)FӱWGX͎͠i9���L��A�*�q��+\���v.$%"P�?�F<��FA�ȍ�����>P�D�[�s���A��ϓ
6r�N��ｓ䙫���;9�!�^-�G��e��GK���Ec9�Q�9��}?B���O���m�L�=�B��NT��hxpgy���3��u���X��R4��� 1�MW���K!����tNU�p�����yE�4~��w�Rn#L��nH
X9�f�'�WR�ş�V�gVv1�I��Fn������/��VS�D̦�$�����$�x&3/��x��lh�/�}�C�_2{�2�"��^?���D�6>+U�6Y��V��A(v�����D���x���*�P�6U��U@ �e� �X(춧�.j��f�/��\c4җx{Y�{�cs ��f5�l�	F���ܪC�k�pf�r95��<�E�SB4�AGX�0*�.��g�$d���A'G:�I!�/Q8'�ԍ&���*���B?�3A�����Z��^<SI��FCg�/x�.P�z,�	�܁��}ݤ�*蔵�a�$@Ɯ#	����)�5��/����t�V�`�5���ȶ�ĵ���T.��Dyȷ.�U"|c�k��E||rF��d��pӼmO�����D��2�f`�@��\U��5�Rg�Ws=X��(}ӎN��}S�����p�֨���"���͝3���і��CW��Q���o_��b�� � dӺ���l����PW< 勝{࠻Nl���}�d������V�*��+@�Ю(�b�g���,�K233g�v17>0A���Y7�@?���ᥩO���#a����c__-�+�M��FH��iY���Bk�2{4h�[L[�~�4 Q���8����W�D��NO�T{�����ܿ���z��`�������;�v�oN� �Z�����̸����l-q�H�I�H�Y��V���cN8����r��S�ayI&�cB#U�'`rߣ��F@#dh<H)����� k���NxR���g@�\@�C�,��HJ���"(�.���}m�[��E�o���Oz�[��+������K2�}�]O�\�W"Z�>y�g����'�U�tV�W��ݿ7R������\MX;��#���j�+ڡ" �>�s��-������D�X�/͊�g��J��+�Th�G�z]��d�*���x�x<k�z ��D=ʿ�J��#X]��	2eL_��-X�=����	Jc��+g�x�R�2N�8-'�f��v���G��Ԏ�M�?7�'�N��PvJ������sW��km������*��-�7� ��k�t��J����{��I��/N �_%b#�1<[:d�޴�6�E��ƨBWoj������S��'�2�Y.���`@���ο&r�@�O��G��%j{i�Y���t��S�f��u���$�$� 6�����٭���/H$~.��[��>�����"�����h�8�3@V��M�+4�	IA�F\guQ)�`��P�!�T9X�]ʓzYw����;:��/��I�c��e*��.K#�	D�s���Qi߸��\���zb��b�@�5���/a�W:q�$t�ۊ��8�����F�a��K��MŊ|/��)�z�J�UZ.�;(�r�'�SI���ϭ	�%�6��ӡ�&���7�u �����������	&��	�?��	��O��u�{���V���o�ͭ₶:�W�쉼���e��հU~m mx#�c�ھ1��\��A�(���[ˁ�����h�D�T��<BO�dL4���m��T�=�p#�U~���#b`�y/�W�#Rh�sD���+�����b��:��"�ZE%j��@V�EA�N�5"f0��ZH�3\�P���>�'l�l[�1�ŏ{u�~`�A��Nh��|s%���s�Y]��Gu&�n��[�~�r�|�W��΄���'����jE����AP�D��wH�s�������]��{��E�_�Wܾ5C*��I�b!�r�~��Yp��4���ο:��BTL`7D�����v�eR,��O ��ǿ��f�Y$���T1�D�����n��L��< �v��œЀD����Z	Ta����*��	��h�����������1�UM���j~ug<!�L��ouο��k;ʉ#��#���s�8��&\�d���-�G�_�yI�����O�����_�,��츦q���[����Y�J���3�\�o��C���f��e9�Gv�
n���X`Q��aq�/�l[.�}(�0�3B�U*[+���;�E��o�)����2cg��K)��o,6ڥ�=�_%���y��-#��-���@i�J�5��4��ϼ�|��7d�����ma4��}ro�$�����?U�-ʊm���3\��R(��m�)�U0W�ӥ�����t-��"�M�l�\VD����လ��׸�k4�"6�
�}�����s]�kɴc�~�eӋ�r22�q�:m�P�Ks��[k?1b��s�����ۺ?譤�2&������\yXN�ͪ���U=G[�����F=�νR#W˞ig/1��T4����wI�@���X!�x��	��re�O8�p;�Mb�wG�3)9`wX��҇�!�Z�#m=���jP;t�a��N���Uɧ$��g!��g�<f�[���ï��e[���苪3��~�bw)�E��r���#�5F����or��w�F�I�4�M¤�_���������=�#��K<V�ڱ)e�.�
��O�N�G�TԱUK�� ����5�.�2��O�Rk�M+��x쾦�%գ~%��E|l�R%K{d	��W7�M���=�w^�d�^����Y�E؆r�2��t���|�J|����>aX0'l����.���Xe����N���GƗ�\(�O�Mj(6l�%��;�~z5���eP���i�����~Nw]��� �d���ێ��O�m��^e�!���h�ǽlC�\u��}����T��/�k�]�������sc��N����A�
a��Mx���u{$A�n}�,2*sЙj斑�_
�?�Q�t�\�1�麐�P�06���w���,�I�o�j.>�F�����}��˽(�|M����Ό�6��z����P��Y�D��S���_��]����q��V�c�7bv��`�$I+�l���d)��E�g�l���l�m�h� ���ɲ�"���?>.�iT�3����Ooxak��F7'��s��� 轢�*��'XU����!U*r<l=�<��˴z)׉�o;LKe�?:��|��-�����L����r�H1z�؛
�����{t_�F9�̎^Po���7����C]�c�L�/�ޢov��|��!�K�C	�wM嗠� �B��Y����bi�c���5(0%XJ��w*�13�����^�ŀ��0��_1x�l�P���½��y�b���YFx��鯻 -��H�I,���}�M'��o\���m��%�9x�ȭ*:�#M�C�i�5���g0:$�<'џ:l�#&��Y؆����rW��W%��e�ɓ�d����Nq�j�Ά�P����l�NL�ꟴpg�5��{�����w�^n$��e��>H�c�������>���z��0j�z6��TV��~v9���?wb1�1�bo���vW����[�(�b�9����5����9���b���?c5a�@��"\=��*�@��[#��/��d�6��nы��d��K�~�*������b���z_���-�)��"��/�@�ͷ�eaؒ1��l��;g�% �=���+�✼�Uk1M誔5�����J�gpo�\����l�*Ÿ'��jx�x�~N�-v/�]��ݠ���Q1PF��T��[�i��*�ڷ���uU7��M���&r�i.>����{�(���D{h�<`�T+���D�^w)�<��2�b��w��1�N�fe��C7S�Mnu�M(���7��5o�K�Ժ�ǉK#}���#��M(G�q��2���$�����Uȫ^�oEĤk'&nu���7���~XՕ��ۚ�"�40�l���jA��	�㋕\;��,��wR��4�_?+��9A��kpbv�2��p^>�~���盐+�S���.�>9-�Zz�9�ng���x���so��(�s0'�0Dch�ʁ������N-%i�$��+a�@�|#�ks$׮����Y
;¦�*4(�^����*c����&h��ikS2A�Zڕ �P�\�u�q�U��Tjͧ��F���p/�N�v�	jU��k����B����C?�	?/yQ@%�M�_�'�g�=|�/%
x�����o֡���E���z��x��iט���]��b���;�bͿ��RQ��Xo���¶�5����]?�V$����('�/Ʈ�L��4���~�����8k���1}J��c�I�Ƀ�(T��14��(S,s�%@n�U�xjm������d1�7"F�Y��o5Qr�$�#"G"[�	"+�8���V��iuH�^�BU
�����]Q?U*J*�H��H����l
S�;��&�V���%KC��%m�+�}��3I7G�iQ��̿s��2b�X�Bpu`лv��<{�x���<�j]j���j�yU?'�	�S��ne ���ܜ`�R¤�=�o!TB!0פ�o�$���kYd��|�F��*�~ � �Ll�N�ѳ�\�L0^�x���M��'��	?Hf���a���䅬#��X��� d�̻GCir��f��m�
��L��X��h�kj����ݱ�(����B=k]\�����hW�]IW9�����91�[�]0�Xs���;P������,�1��*����������'%X��#�0_��dw�Yh���׉~)�΅�S��/0WVG�:x4p�z���.̮���ֱϥ?�� �;�G�.c�;a2$���Nv�DJ��eD�._�<t�El�=�;�����$��#J�G~/���@��em�?Z��R���Ǆb��7�K	Ő�q��ei�f%�v��=����-VoO9$3[�C��`��Öp!�}7̿}�y��ׯ���9.eu���f�'�*߇�S�P<���6�V����<��Thڈ��]H���;��X��J����^���>I��ɲ�Ne��>b3�:g��srdl�@��@�@��@���E�=�vg��N��&������>�5���K{�\20�kK�5�����9�r7/�&��8���}�S��Zay;i����P,���AN|��[ JZ�N%*Ҋ��~b�5��8��D�����-��&�K�t؅CLRvf�L7��Ok��ظ'�3$@I���Cy(����A�,͘��`��0W��R�]��S�qus'�Rj9)T������Lsj�o__0e�*'&_�,�oƧ�-���Q�p��s��Uŝ�g徭���@��>�;���z%K�Qm5������!��7�>_����^ߩh�+ҫ���$�#��w�4a��3�g�/f��T����ϙ��@�o�;^�pn؞�|���G�C9(�����pcZ'$r�S�����MV��w;���>���},�F��T0�f���Y>6�*�B�o���{��!�'L�F'S����	
t�<�ҟ���fހLlGt���lE��@8�µ��]�3��c�� CO�.�N�Q�cT�%��g�h�E]�2��Л�Sz���M�쌋�|�}���z��3.���8q��RQ\��b�ӹ ����\Y5K���0� U��Gh��sm��+�rO�;�����5+H� CY��S��}���~
>s�?D�'D�`��a����O�J�*	�-��T�镀y��i��ۗ$	UND��;��ʽU����a��$)�^6	G�R)������)�D��="ڽ�y��Q_�'?�Y?�sj��;��lۜm�/� ��$GF]��4:�7G��h�m>���tʝ�sv�ً�qG؜�5�#}�x����U*�� ɿ��%3���HE�"ym�f�.�c�"w��Xg�[V����μ�C;ɣ��u��� }0��|V���@��Q�?�S.�Ύ}�^�6�;88(޿���f[�wX"�e�}���,| !;�z��	������"�<ۭ_`�ғ��Y]�~���, �������2���O���H�J�6�+������|��i>o�+C@�jd�τ��cs�VT�n�~�j�<&�,Nc�U� ��y�;\�Ȭ�=�s{2n�g1��S��~��X�K^���У-̽�d�Pz㳑��&���� "�=�(��PY�F�P�3}~�cb{�Y�	���"�w$��NSf���0�Dn�-�����س� �m˸+�?��Ky�F�Ps�_�}x�'-�ol
�'�ƭ����P�-��KJ?W�t�s�Ε-�f�9D?��{~q��	Ք}�}������\�d�ؑg����ͤ���\��E��sQ/@�;�����
�'��q��c��`e��4�0k��nn�׻��h��HN�6Ǒ�Le���#*t���/b�m�eέqeӭ�`�Z+}��-��X\��� >ͧP�,e�m��8�TEI��e�f��j_�����]�cY�� ��;����ur���3J*�E�n����k>��` &�w �Ċ\-�㲻��/�Q
1�(������DƖ���C'G�_�Н�;B@e(�/��e����͢�_�H�0EdFk5l�U�	�Q7oS:��a���D��PvB��l _��{�ni|��Ȍ�8z+������v��?%�����"��i�A�m���[��������v��u�%��E��鬻���5�~o��K���	�s����`_�R�	�		�y�@0�l�wU��m�v�B�3�
����yyE@+hD��B;M텁��=_ov����C�οb?9�LLP��u��ו�^��ܴ������2k�C��پ��=Jl��ޯ�3W����rs�
g���T?x�9
�W�t�9���b�1�K1����fY�2u�@���:���î�N��.��6�#l2|V��i�O���$�d�\�9*Q�ݢ������a��ϥk��&X%2Z>�C�K|�@_3^��e����_�~�ld��L����~��7=�P�ȃ^�9�[h�|(-q@xt�D�����n�F�2��q%R?H��|Ԥ����TyZN�a=���@�$�C훝w�,�quz��%{�NO�����3�T���(i=k� �:,Վ���=�:Z֥�ݦ��?�]6�4���Zu�	��w�R�|�~�I�5�w�O��F]�iq�f�`�n�{�N�e���:#�E�:�w�g˯���xnƟT��Y��Fp�K��ܜ�;��n�jPX$�� ۞(��E�8�������i��A��sA���G.t?r{�`P6w�����]	Mc|-��q��E�����g1�6��yr*5�-1��w��f?�(�(��D�sC�>f�+�
}�ﭛ7%S�&��
�m�j켪	ڈ���smT�7�y��t>�l�+P[<ݤ�����r�(d����U��/Z;[��� �������f�Koc�7j��C�P�݇�L�������]k�ͪ�s��v������?�����*�J�Y�(�gk�����Q�n|�1���AM-l��_����f(� gV��xu��>�6=`߫'�PОFG$!��%��N�X������Y9�@l�s��Nh�ݾ*�T�h�k�K|q���Y��_���8~���
kpxR��B�m������3��F��ݰSfC�]!���|�
R;wAx��_�>��6G;7�lh�n<�	�ʒh�-��g�����X�n���m�=?��ӂU<^[����#3IrN�1������.�ڡ(�~���_)�E�e5��dTO�Ҟ�＞�9�^�ԅ�M�5���Jij�\ṩpz���is�]<DG��>9B��4�{�e�mysD^G������y�[uq�+���*�N��`ܓl/a�pC��ևg8I���R�iX��@���� O5��,HP�$|#ٛ�"���b0��ZLP���� �.�QI���N��0��NRmzO������$�R����ɓ�*��G/N:ZY.5�+m-R-r�!������ڹ��-!t��I⏯�������T�:e��r��^�VSDk��x˼ts�a���Ĵ8�]�K	�M�*�P��P�C��΀��-��d���M��$N/d�;�=�M��յ�S?uv��tp�P��t�_G��~�v���m!�ak�^�����+�v��t�L.
˭�Nܮ�'��?XF�-�\�,DxKd3��/{Яt�ǆT��B�Eט!��@��^k?Ώ���9@�����Z`�}6ܭ�&�����p����:��A	��;U�7u,�}@��p�����
c�(ڂ���	��-NO�-�eMj}D<H�A2R-m��.��YA������u/��o���9�N_��%0��0�:�W��k�V�M_�i�Ћ�^PGq����e�~�r%�g*+�Đ ����>�4��!Uz��3��8���� �Chm���hdndn'ܜgaL�?�d���J�刺��J(� cR�����,s��nު�H�V)F�aM��&��m2e̬��O�-�2㷙�xs9+��j�
�o`7*�U��!O�+s���=���9�>bq#̼�W���8�@]\+�KtV�h�{8/��ǔS8E�gms�zi8������t�-Ѥ��(�{�Ye�& �-��2A��ث>H���sD���1���3oEWi�1b�E7HȨB��}�lx?_��WpPl���Z�z���Us�*�,��r�,�[7}���hp,�5��
D#q�/Fr}9^�>0*�b��#�)��[UKٔ���Ybں�2������+��Wg�D�Q&���n���{	�P�����+:ϣ\$dRQԕ �f���,$���3]fk�Pi~7mG��4H)Kv��m�YF�=��SS9��|���̳$LQ�RŠf$�#i3q�q��'��N��E�l�(;і��|�^h��\ǟ�4s���J9�<��f7c��( Ҙ�L���
����[��� ��=?� U�=�]oGv�DqC*<�QBXJ��uu�ce��sA�č�#\�=$V�����*�G��%�� �ι<_G�"��%kmn/>I�������������.����Q��v��RS��X�ty���sN!|�w�b�z���Bjہm1���ZA�&y���e7��e�X6j�8L�}��l��m�7��&��%���ͥ �Y���{�,Km��-f�`��Xy������Vn����lx���9�7�2.�<"(5E��N��e�#G���T��::��� EP�����Nk��u�c9y�J�z��*M�_'�(8Q[�t��6�7
1Zr��v~�Ѕ9�L�߭q��<eKW���p���0�m�����qvHz�R�./�yR���9���&2����mln��6����N�sx��2��j\�#����V�8㻚�y����E�g�V?�YƮ �K��^� ev�%���/"��c�IR�f�HC8���j���`��U�8�_����z���v�0�f�y9����CQ�$/�!�R���� ���7��b��C5���:�=�"���ͺR>2��$�s	��V�t|�~�-��WN)������#�OW�Gphk�d�u�1rٰ������A�z�S�*�Z����Eoh��y5���*Z���Ї�|���N1``�g�9��1��L]��r���N�C/F%��>9�Ŗ�l�W���y�=* ����H����{I�O$�$#1��_
�{�L�q�e�����L�% r�rt.�@*#=7�B3�J�>���"�s��Dϸ��Q_I]���.<��L�����ܠ���-�j��m�E+)���BWzS�|� ��媒M�%q錸�`X_����ː{Լ��J/�D�m�gaPJ[�|�4{��nnr[��'�*B������b��GF(�oc<vբ���J��ͧ
�~��|����}�Ev ��bC����¯e�����:Yw��X���F.D����(^�a���Pًi=����W^%���`'��˾���>_/��	����"�l��%y�k��k��*ߐOr��|i���ׇJތ�8�Uz�N�eX�I��
��P���LO�z-���ZQ:U0(AF��'�6�`���z��o��\FE�Hb&�^\H���U'�b}ߟk7Ql�~�>�X	�������W�<}⵷�n��z%pz���}�$�EkN�ߚ���>|rf16uDsX��f~�Aΰԥ�b���7�����+
܈gw7z�PaG��Q/ة|S7�+}�֊� E)�"�ĥ�>���>~w�HW�8���<���؀(�(���ĳ J!"���lm>��.��K�~�d^����}F,(qE.�B𾥎���j�s|��Z_I��s/���YL�U�0{uH��a;@J%�aY��$��+#% �:%���(�7*��%q��8�*���#v� �S�]S�-gv��d�xw(�7vۆ	0=�?	H`�)��'m]%>�e���IRg�f�W���w4�)!�8l����~)[�0�t+���}PC���h4��s�=H�]�u#�۲�xTT�����!�;��*��=��/v�64pՊ�H�oX�<����y�:}�＄~*����,.����#$_�P��[]��74x�e������ޡ��p�Pr�͂�����5����C��I�Q̇E%��0�AY��yz��i�)��+݇c}� �T��k}�j�	��_N�(ٙ�)5q��W]`Tꔜå��?��p��x��axB�q�m����eevE�cJ�~z݉k4�f1�,R���MZ�����`�|��	��\�0�s>��}�cx�u�%�����aaz���W�����t?(�"��e��J��N�s��}В!b� +�-�=�t�ЏU����R�֙��'�ݱ��G�z��{��]���TF�>fV�N�����i���'��&H|$�%'n���K�7�+V��k��AKJJb�>`��K��*)SyZ���5D�/jpK|�o����?ww�������FT���k����%�g��[�Ж�0�i
�>��m���q��3%VF��H:��ݥRW��ntQ&\$��20�����>��L}X�@��8s��E�۬����Tj�,�ድT�8��pĠS�xo�(Ҳ�B�-5fM�줝������0��{�;}�k����Q�>�6�D�4y(�A�����cz�������N-j�?#�L����"�)/�;�Ԓ�?^O�A�F�Z-d�V�E��h���Ou�[$P+rŲ�v�655N� �H�P�YMA9º�ʸ9��q�����-���	T���_s����xa�n���z�ա�5�o�����ɡ�`���j��{UM����x��k�s�ߨ�i�@��?X�����`�d�!�I�ŖmN*oM�3gK,�
�E{:|@�a'��,�S�?!�*c�����$��!�������/�	�@���ޯH�����%��;i�g�d7�K}v�L�a���87�� ;}�*��l�����Cv��]M������ت�?T�����wC�\�J���f��KC�
���MY���t4F,����=Y�4���i��%��Q惧M�%!t���S~�����Xmv�Á�7���\B�E+�'���U%_�~��B�`�T#�(4��\��8Z�Wɳ�� ny�E��p]Ͱ49�@�p�E3ApҮ�-����%3����������4��[ϵ:�|��Z[<��)��(y��W
�S�T�W畝���&�n�9��z����m����p���v�������v:�Fʭ�������Y0"��$���T�_~U0�z"{Gwc;碚�t�ȗ�/��r��ث
��5���,m���ZWr�_��D����~>�-j�ؐ�Ө��	��'��PyՓ���<��xj��6�QB=���n�A��z0Հ]L��e?R�V�y�p�\�у��	{LKm�������V-�1�6��:�Ǻ��Hj��f��-���s�5��2�3�?���vk���s��g=l�5G3|���lW�B0G��P{�G��Ыm�_:a�ܦ�ߍ����)�K���g""�Y"BeR�Jٙ���}�!5ʖu"�(ْ#D�#;3#Yg�1����z������O�{����|�=�h@ɘ?�Q|��n��*��ĕ��w*ZNS`����::�Z�`&�fϘ䞌GK��@׹��%a��l�WY5�~XI�I��(��;��x(�T`�5�S�����Z�O�K�|R�^�É��q����
�-c����,i���QJ����O��B��_��5?^��T� ��w��?����5y�p���!���C�s�z�<��{ҧg���7X=o�/V�xs�����t��R�+"'[޹�XlL>�0� /�sn�y!�J��ٻ�4�}}���%�/^�a����|�_�;��+:u���������[����%�shlO���F���[��˖�d����3�̮G$�_��y u&"�⬃i�'\sE�����<Y�K/�
;X.�+7T�0bE��|�mؖ>w�1ӭ��m�o��Z��]�%�%S�	��{�^F�DbG���Ql�mN�k[��n��;�B�ofG��| ��T��c1I���W+����}���IfC 9�x��S��/9κ�oԪf�fd
˱��
X��Ň"�w����?�o+�?M��L�Yv�S� �؇
L�Ja���j<)��f����	��h,�����?(e`��Q���1\�,%��å������"KA�M�쥃���Zs垹�u�ep�	����Qi�ق��9&-��t�r�by�A�e�{��C�(Y���O�0��Z\K��,/,&��d~�d�k,���1ߔ��LY�J%�X7�7l}�"�[��(��G$4�ƒ{&=Gb��`����F��O�q=6zҝ&�^0K�P��|'�@�oIU��3�y��SW�Rz>��lJ���) W�O��0B�gaQ�'�L]gݱ���x�ѓ�n�W��������>�)���GqCE*t�?����Ε�Z��L��!{(짪}\c~�Ş8 ê��P�w�jw�p_��O��u�@��ӹƼ��|�\������뚍����$�p�|��Ɨ�� ����E���n��o1�th�7V!���,O^B{�9����*��E�*L+.�}�)NT�f����i���3e������D�Ϋð��&/{-I�d������2c��#AW/D�� �HzP=+�ve[[[��M��Y-���K���$�R�1���L
_�q�Y��`-8���Į��d���@�~Aǰӡ���x%,��]����T8IݺLθ(_������$���E�g�ޓ����+����(�h3������2�HXs����N��Njx�k߻z���E������:Xb d�.�gkM��3�v-VxƂ�g�4롬K��vx�͙�V$C���v�v���� r �c,/�ǟٮ���a�%k���{��ŗ�#��c.t�U��z�>9�� s:�a�j��E�ڶ>� #*pmuQ�w��r5�!Y�s���c�.�*����%�2�����Z�K�Jt����ޝ�N~���'ڭ���
b���!�9�o�PF�Ȗ�N��V�jS�bt'�˖��y���D~]̸��C��d�O�PxZd�N��sGft_���"����ڐc����R�EY�鵊o����ʻ�[Y��J/弅Iz��*��cw�c��CB�ֳ����3�֋`�ʅ��{{�I�Jƹs�<�9��n�|+�FG��y��v�����~W�e�u�n�p��*�<��i�M���#_�@?�[��)���_�2�@�AD�~%�q؂�3.!;��?L<��T��Me���i ��V:�����7��
Qj9]��\����w�:��s�X·7*��͔�������E³/),���8TI\���Y�	��@���,�p
�J����?<�E��?�I����	4�Q��ȯF�.U�rx�����/:���u���G�*b2��
��_��^��`_@��)��݆�y -.E�<%!K��dZ��?SlTZ�G+h-h�1z���E�1ʵ80/��<���V�BC��J$���GNCp�N�Eab���B�Ӆ���	��.���ýE�����pp�F8����5O\���󀕾4=2�B���J��3<�a�Ǯ�I���7��!d�h����X��olf/����"�<�bw�Et,���@��H���k\�L�x=C1ȩ0���p�>۸���lG��Fc`�K>��@Y�e��U�~{�l<�yyC�m���jw�D_���۫kR3��w��=#�CP�~�6d\���C/�7/�]>�`t��t���x��+I������Z?�7쒡�Q4n�`���R'~e��.�3m�EA��Mu�M�?�ľ�/�؅���Q|��A��/;���ݜebnC�V�4Ю�_OO�}�z��-.r��mW2��?�$}����-,��ǾeW����(��*=��>�BkͲ�ĵQQX���fO�=�檭��Kk� ����N��/~���親Rr�R7Ý[R6}Pܓ#|�k�lR�E;���~d��$�$n_�V�:v��YZLOawލ���G�T[��xTz�4O�g�#'�!ъ�-��?*e���Tl厯(������)|�f��u~eЖ�K�w�_�*a�D��1h�Xk@��cva�mZ�d�wK:�<��㯌]��/��+�wND��}ey���k���˿- b�ۭ:Q�+R�|�B���ƒ�W�]��9f}�n�U�"D��u�Y/�x��d�~�	P�gG���[�,K����̌g�$'���7���[���Շ!�z�0gM���#V�{���������Ô�MI�����nK^8hZ����r4�0����I�T��7�S�*s�=���^V��p/�P`G*<��m>1UF�Sz�>�pU1J���]�k�h�Б�pNm��Xj�`K���zα|`�W ��oa�\m���k��G����0��6�`�K�Y��uo3E#F�yJbb�=��%����UX� c���ʭ-_�|ݎ�l�k�����V/�K���4ٓ`�Wcy��M��&� Q�TU��\�}6 ����ڍ��$c���a������k���Q�o��m&�U7�}[�{��Jw�q�j	�4�9#u� �z?Y�<���nG�X��`�U�9��&�����E*��[�!��������nsB���ި��5���=�b��A�
��:�ur�f)�����X�S��'���H�� �-����VPK(d��`��Vi�{�ns&+��^��^�����镳���y1��>�o��W�~I�ŠȥG��C��	��wD�>O֞+�Ô��>�.jr�=��t6WjUڬ^�΂J��T��Y��^�^�]e���֨ADr4ˆ�G��� ���:zM��}EU\m+�WP\�ɯ4s���e]�\	� (�`+]+as�j���9���JP�<f�ԥ��;�:��+j�yn7.K_��c�D�ô��ع6'�����/�W��m4�/3�ڄ��	԰&��fZh��|�W ?���I�=�Λ�*��4L߫p�A0b�Ƥu[��͂�%@,`��3�����q�{�0Dߚ!=��QO4n�ݍ�>���m��D��$�C��v��g�Ä���p	1U��]�7��W+&�����B{�P����fI�� F"y�A�
��bW���;[ݨN	��$�>�v�� �%�˗D��E�z���	;h��* �y�Ɛ���.]��)��-/�ڶL�abh09�n���� �Ly�]�uԵ���|sR��P�ޔ�I"�����j.���V����?:	�q&p��A�4-}��L^���y��$���<��g0;���=��)���ޓ^�yP��ط-&켵��}�%睡��z�g>��i��Uz���;9��Nxi�[�����З�� ί4 ��b��6'��J������1��g�l0��.ǽ6�:�_��@���ez���.��57�}���Д��fHv��GeZ�ԏ���q�'�]0E��L˺��+��{q�"�f�I��K�|�4#vf��Hm�=��u�󨡖�r�p|�?�*��sºM3�O��&��U��#��R��L��������?x��)p�N�	[JW�b�L?<�l��C;;�r��������(�/s��+Ն7�]�u�]zz#�g�b����1?c>F:�i��`�l�ߕdv�e��4Q�>��F�f�ǌ�eF�C5�Wa�v� �TH\���͂��,蟝��\�i�CCڠ�E�u��{��
n��j�ih��s w�
��.���!3�1D?5�)�x�(����]������2�kAѪ�Lp�_]T���� �#���夒��ӞsR{�+L?����G�T�"aI���PQ; �zG ��8�/?�>����4;����S��4IAB��⮮�]��GՅ+~�]2�?������Z��,E�c����
���� ��Ժ$m��� X�pp�UV
�x�a>���
}��Ν��.9��ث��x�اAC�]�~��)~}����-���J���{����kH���A�'@ɫ=�(�D��A��ʝ��aR"xY�O���(y�E���}{�5ۃ�Q��Ĺ!���'�P6����@�+f�%V,dc��5	�:k2�4@�識��2s�>�����B�U�t!�|��F��K���C�G��&��N�_@R�f��GF�RO�G�|�\KNԺ�W}�W��B�9�s�7Ltuu���i?qB��є0�v7d'����x��{�P6�*�S�\h�����A��
�#;��V?`�����5&m������R��~E��'�o<� ]�w�3���2'�t23����n#���D��>��Ѱ�=B6���dt��gU�Q>צ�HBp��]�'K����ϏW0z�es��0uG Mߕ�	��HC:�ZU>����)���y?��\���d
�����/������E���L��卿<9��^�1�_��¾��T2/m�����q!
�|�e�nЙw���~�ўC�ұ,�X����c��sEBѧ�����we��W&�'�ٿ6�,���7{�����s:~��e���b�H�b���4�n\�,V�-����]�I-�}�m9Z�?T���D����qG�4�~&�?��-%S����>?L!ZD�$A�]�u��!1�����c[Ɯ�/��zg3YKsɜ���Tk/$y��
9po$~�)�]�t����x1�(���R�����s�ԄP�3݉�
�#�{(�)'$��2*Z�V�i1d�����5�sV&a�F����2��R��>���m�6I@����TL<.��(��$���uJ<pŐ(Tc(���D����+����t��{�4w3�y�[����c�LM�	�n���~��x�<�hr�Xޛ;�
�yp�	rz�Hv�7xy��l��f[!��p^
`я��}�����z�r�8XTT��\|lx�>�!:Ŏ�#��J�N*�F?�bP����Y�v�0�\�Z�]�2'3ܮ
:�\m;���f���6V�|MO:q:�
~:��*�a����#&��u���G�x�k�����EWѶ�R�]y����-N�!��v�p{A��!eMJ��N!᧶����-3����1�P\U\�}�7�'P�TT�j���h�rG���Ў���^��j,s��
>�7@=�w�>���2yk�\%�'��� �v��Q�fϪd��C�mf�1���>�����
�A�拢L���C�k�f&Nv�j"��;���g��7�,)MZ�:M��l��'��P�{ �ȇ�p!�r�������8�=�"�?�BΛu��\�8h�Y���\$�����G鯊	����Tz䲥���/"����V �����]'�nG��Oy��u�� �d�:��!�az�߶�6y5G��w%���f>4|ËmG?9�Q`G�A^�Av�ɼǉ\�=q�˜��'[Y���Iu��v�����]�/q?1���r+ �y����SV F� p�s�jDb��a��x�I��g d���%�격�{�_��]l��p�V���=\�_TM�M7un��)������*��7�ƹ�A�����%�h�/�D*I<���>�l�\�73^"gD�-s�ƸТ�A�!��0�[��QON��r@ve�$K�]��o���sQ��O]�p��+ ��N^�,��q���̜�O���
rOC��8����Ah�/]"Y�@�7��9����/�X �T�4�D��	��/1w���v5|�8� tiU}:9����T�H���$��6�c��:����2�����͎��Ds���e,J�W�f�E�J�u�K����a��w�ׯ��|��E>���֑|(��5��b�tT-JL�����^�gW�\�����U��d���t��V����ߴ�%�9պ��lڸ"���� �"�H�>hay@�dcƠ/]���qQ<n���us���ۭE3bB>g�\�� G�̕�{�x����y|��)� �=�'B'����k��1��R◡�������w,T�(�#"���gh����R�\jD�HʋXe�����������i�
���˪T��xpJKw ͵1�p�1���Q����fo5W��~0��x;�+��|~x�m�$�'US��Tp7�$��~�����X�����>8q����E��sИ6�!�>��ɧk
���`ߞ�%�����ޏ�#��
���8�q��vZJng}�9t&�Z��G�{\�9������#n}�;��J��Č	��癆n�%����Iy}w[|�N]b�tCm|ץU)�b}�x|O���G��ǟ��4�Z
i��0�=o�3}z�
�ΌV%��t�x_)�N�H!��[4�����?���W	�t�A�m�'�&��U��8=/q �d�����N���78�_:�����C����ͅ���ى�ma�Yg��T%OL�h�Z���d ��7R�M��$�����*Ҡ�����ڈ���E-1�xSXގp-��2���v�m�1� �S��a�(K
]`�-�}�E���*����QG$!N5v��vz�)�b>�q����18;���אe^�q]7ׯۥ�tv��h�U�$�=�E�8| ���!���_�ͮ�9�����-��w��$)H������.{j4�],E�'�"��;7�DP�M+5��gq��;r������A�mT���3��K`��q���F���
���V�i�?����l/��hT��M���Ă�L�R���L�("��J�5�%����-p[6�3^�l��ѣ,�r$v�����W��}����D�;4��]��[#E�nJN�&X�B��Fl�u��:�=��Ks����^��[�Z�m
�Yz��̯	`���W�j��{?�Pi�H���$ㅇh�6����8�..��n��^Ҭ�x�som8�����S�� 4�tcp�P�2�U������Ά������Tx�l]�"纝PQ�U�I�M|g���U|���}jhY졈�Q�R9vW��^'�W����H���S���B���S��(!�Ȕ��W2�]Q�� [͗,r6Qi�j����wg���
���R<��v(��[�Y�H4֘����5���1:5�d#|��:�+�O3�&���O��S�[����sHUrW���*6�i��ɹ������ʡ�k� ���&(6�q���GO�8��U�u=��X��~S���q�?��O���❴
;��m�ac����̿���a����41v.�P�48}@����\��F�=7�/E_r��1|sQ�a.�m��n[�k�K��g�z���|Z>![rq�>+���N�k�3b��B����-r*g�]�,<�܀�J��BX*��m(�?���OZjYvR����x�ΰ/ J�o|B�̧z������6�?�m��)f��r�\��w����L٬��Ƅ���%d۴>+��g��u/f$y��2���"�R�����C�Ї�O��v����^M��TGV�Z���k§���^(u{7s5��'�a�n����E�zG)F�O;�<uI|f4�� z7g�$�r�݉ʫ��7�=�;�۱�� �$�6��hss^�x9T�;��ᔄ��ѕ2�qC�Y��;}D�wǓJs������B���}H�)IY%)����K9�Jy�����A��a��@�l���i��JK�"�9�Qr�eyW���RR���呯��7����}jYk]XL�8��Vn�gCHyx���E��뵓��n�ā�e2U8W��d�2�����	d�M��j��iW�W~��֢CS 6$��gA��ЯʒE����3
5�7�l�-v��>CSXfX��f6/��,L~���e�ص���b�����3�[E�D�#�9ky]��i]���9����{i�lV��g9Q'��Wa/�`�W�6a���	�O��=%W�o���QӃ[2�J \�o6��[�N�_;C;�6xߎSν3����V����ñ����z���L�L[��"��ɢ6�����l'�����j �frn8���$
�^]4��Ua5��T,4�toO���1�ޒ�h%�����ר�Y�;k�xb�J��ͱ�/��lZ�--L�s2�{�WGD�Oέ������lT��`
��sܞ4��*����U����^�*���
�zZ��Aݖ�I�:);��X|#ݕe��}�c[�A�r����C���4�?���*�L�P(`RW�t��sA�?�%����VW����]P��ˊ�vWص�l�}-I?�J�n�Co����i�쨲�"�����O]�艏4Q�w�+M�󸐉<��}S��M*��ג�����[����vm�S��;jŁ6G�����h�>��WX�p�V;$4������T��6tUl����R:!L)�O�_��8v~T���T�I/.��3��N�w���((�^�85 t�6�L���=��@���|Z�?���=i�l�,Y��_[�?JIU�Æ�J�����tZz�-�V���1V�S���V��m	�~S�yj-wğv]�N^v��)�_��1��L������A=o�L3=��;&�)��U�H�A�~�e��P��&�̥��w��GØ�Gb	�����]Fr� �eK^�����v�U�mu��e�:�".\>/����E��^9�X�t�i� �(�=���v\(��#`���\(�����cY�n�T�uR;����yW·������:_�6JU�7��w-Q��eV�>W&��sǹF�R�zltu^�c�L?�۪LR�6����ø�V�Vmq�!緈f 4HC�V��Ш<w�*���:�zH�e�=ٖ�&�V�o�{��2do߈��<�6�+�*엩���հlь����x2��#�G���f��d� s�HR�w���R,��M5�u!���KՖ�M��},Et���l�'g7I�ѽ@l��b?}�/.��j��|q�0YurM�{��:�f�Ϲ����>�gw�*�9�0�02.1���n���F�X�@��	ӽ�4�x��EC�=�)a��~�n�?|�����\�-��`4���{��`=*��b���0�� -L?���۲
����C�Tp�@�����<SErc�]&,����R�k�Vz.��<�����*w�
�=��>���Vm��4����� hExt;�t������yH�Z�߇�d?mO�����a���G��\�0	�	�j+P-FjmC�F�8D�=1��m�������ESSΆ&�;>�Ҽ���\e��<��/z�kW���NT�F�U�(b��S����������	J/���)�Zk�sc
��������T��Ӧ�����@v�(N�����"Q�]-�}�h-v�y��	<O�%��o}
���@ݶ7�Kްy��l^�s�����K��=b��qM&�r7bE}56jD���$s�uD�ȧW��5�5d�]�\�[�ɸO�[�>BfG�<����{�dg����;��ww c{q�FF�Cʯ��cÞ���4x�o��r,�B�����XQ��]Q�lo���9�T'����.���'X}۬�$Ɖ�p��ĎJ�\P�7��:�z�$���gQg�E:�UT�(���|��X�w�E��o?��P�m8�E\|?D���9���?�p�v8��M� �k� ����/�N�),�"]�ȥ;6;fyś[r��I(�탌��s��g>�@�>���|�s�}��
��'e9T��� rP��j@(�	�ؠ�����& m�A����{����C�H��4^O�7�c���3����N:7�P�h ������D�DE�1@L�>\[b�|��d���m̀���mS���i9�@m�è ��-N\���e�@�����s��)h��Y7p���]�28��n]��M+P���|ξ�{�!�b���h��A'C�����[D�`=L=�15��|W�Y.�P�rO���d�bl�i�]�C7)ˌƫ���	P� � ��mJ���)Ѝ�`�ԩC���뻘��&}E��FV��c��R�m' c 4^F(��ʞA���R��Ԟm�p��Akd�#*Ǻ1�+P,y���������]���(d��)���E�d���d�� ʺ�rT����k\�J�g��`�̭�����<_:�S��筐`Ԡ��,�S5wR�X}����Wl��<��qS77�[���O��:��L�8 G_8>Z��Ym�jG�]�VpS%��,Gݦn��f�\��Y�݅|�	�զ(�OW��d)�ݰ�_�*+9S�n�,d��P��v�����LJ�K�ߩ�\�]e�;�= W!+���
-�玠���/^�������9�W��n����.zj�6��۞�M�ҎN(B�/-�w:N����R:��颎r@RI�l:�x�>�k��Q��|��}�E�����X�j�P7�mV)ˏ]l.3�7��|�yB&��F(B٣,E�9�m�;G��@�g��D;�٥����U�g�wؗ"�(=���(:@�6OO[U�0��U=��Ο��5W�ǒ�I�`�����,|��^�����P�&y \� Ŭ�v�츺s��Maz7�U�w݀S�P����� ��gT��P`	RcP��Ciex�Ɋ	q�y�x�pmn��|������A�A��34�J�S�"T+�Ys����b�ғ��e:�b[��M���P�j���~��Tg�W�8�ސ��k��p���ԴOk>/:L�	-v���#~j�����0ӏR�ڷ�j�R�T�\�6!�;����\��S��2@L��J*7���.��,����I2Ll��'�l��,Q.��d�v���c��8Ϧx�!��������j�K��F�5�e|�6�k���`
w8Զ�hU|�y9��ܯKN���@���^�F�R�W����ƱC�]�O@�)a����>
�*�*6u�V� ȾI@P�8.�
	-U���nVz	�,\�uK��RU�7��p���Ɗng��צ�hں�����'�Q:�o��	N�u5���s�s�����f��[��OW���;��.��
�{������ Z�Î���#�R59/�ގ*Ao�s�`u�S��Tx*�_:a� �oפ�ܰ5��*������e�j;/T��Uh;��x�c|�S�K����M�FBQi�oK�i%������?�~�m���]���-T�g~�?�d��Yv����)�aoG�_BR��f�*��͠�G��D�f���,�2��!%��yvopQ�sqP@�pͺ�)Fg���kf�H�s���P`Z�;�{�ߜ���:[&&(c��Z��:ږ"�P���'7���a�Ql��<����(���6��n���c ?e�����J��^v�S����M>����L��mJ� S��|�Ț�QW��mR��������r��]*��.�����3��,�ۛ�_.���O9�%s����eE��^̨����9:��r�Y/������-X�Bs�U�I���H��ky]ʍ�ù��q�0	g�c�U���,�������T�i+�S���nqM㘝�Z�����n�c��?�{�ͩ�w�PK   �-Z�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   9�-ZG��{p5  k5  /   images/a528d487-389d-409b-9452-c3cc4275f339.pngk5�ʉPNG

   IHDR   d   K   �"�   	pHYs  \F  \F�CA  5IDATx��}�T������7��{�+
XQ{�-�E@P���Ė/��b�_���Dc��Hs�eY��}wvfg�����۝]v��/>w���=��{���i���6�;>�/>3##t޸�b����RP\$vs9����r�$���Tjjk%��f���{��3�/��������S���?���y�~n����_��i��+ ��q#Gɤ�c��z������n��
ās��B�.��|�y�l��7���x
��=8���rH} �����ؐB�w��5���H\w�<��sȺ�ch����u�z�~�/�3��O����v������y�N��A�x�pH-P�D$� 4w ��|RB��$%�À���-)���[��6�GHDl�����4I����a��e8�X���c���PS^�4���$���RVY!1�/::F�K����Iޯ�T���� ^�W*k�%!!Q"q�υ� ���������S]%��&��1>[W��j�>�q1R z�Dy�����L�b���B\ ��L���qDFDHUe%4�8��QQ��y�`�u�:ID?NH���b 	�$&����r��J�!���w��--!�����G�{�<t�]�1�T��wk�H��\�)y�@�`�D��C�����_���"��@�ڮd8�O��;���!'�($(#G��Z���vJ߾}u��@�ѣGe�xS\�۷_RRRp�J	���C�>%��GP�G� ���s���� L���29|���C�<pࠞOE?��^�g�����qOii�d�=����)^�)���3���r,/O���d̘1���xw�n�@d�R^V.�q��i?�g��J��~�*q	q6����p�(�Ξq�\0~"�Wd��|���="nt�V�����k�>u��_)��TT�uÑ��������%���_j��c��x<�!�w��I:v� �v��2l�0�lRa*3�"2�о}����O�7v��O@:�o/�ڶU���  .���A�v?��0�����x�-�a�>㶞I���ݫg�Z#ǌb"�n��}d�icދ~����9�ݏ��v��m"Z� �W������j�5V��*���ђZlhmp��J~��0��������{� ��dFG��.����/d�6OJK�i�UT��u:<�����Q��^����F��A��q�h?PZ@p��C?u�q;#���@��C�).����7�	���ϸ�g�ws�^���M�{]�n�a���~"=��|������e������[�}�r�M�*�t�t���kj����3�����(�H5-p�98>	?�@k�G^qU��ֱ3��#���.�;i_y���� I.�z�w� ����]����qI�$B��@���Od �z����h�ܡ�^����ݻ�$�:����s0�=�����l7�����C�˞�U�����ۤ�7t�9q�}䈴Kk#�z��Ͽ���!���D�-�i��&� :w��)��5��1w*zB�g���
A7A���������B�zI���t��}��z�t�p�ā-�vz	�oڶUv��g"�ź`��^߳[wi�����zo��t%��ݻ�8H��=�s�T�qP�W4�Bc���@?1P�0���y:�� u�a �b�DP~a�rX��)+/SĽ;vfI%t ���
�K��A��B(��SJ��BiY�Z��e���s�~4�"��'��o"���@8O��u��0r�0)*.�����IB$t��Q���/�h�,�*��{ 'ʦ�ا�E�ܳ�!N�9�]�,�G-8���t�3����B��q��P�/���}���^(Or(��JEU��Ie�k�^��y��}��^-�n�J���y�3/�1�)�u||�k�o~'����@��P��STR��79�c�v �B}�c����5��!T��~�w��,��⩪�8H�\����P1�9'��{������=�ˡ�i�8x�|\\�w�{�!pU�H�@��EEE��)�H��̃�4�r�2"Ώg�?L`��X�x^'e��1܂xm�'���P��~����܅�y�D�!�v����C� x� Q�i������|y�_I: �����m� !* #i���hN�ᆞ�bl�|~7t�ރ�Z�����Ln! �X�t9��=�-�ٴh��28 �@���w���0�����F���M�h��[�� �vh�N�~7�E8u��E���NwX�%���W�kG��~P���q�����%��b�d��9�DK �خ��� �d|g3Jl��F�VM��︗J���ԭ�- �ɛ���↭clMq�->9Vy?�$�`0��ܰ)�fvH 'A����2��Ҡ��$�(�/hͫ��; {'�R�����p���ɕ8tZ��k�GX�/���>���_u�@����jL(�9냪�@0�,ME�&��u2���!L��S�Q�xN����m  'AMs��d� W����q�DB������yd��*�7oެQ�O�KK�կ/�w�j�S�����eњUP��}��N�xrGYE�ιE�\]�O�o��F��P�p`� F=�9PS�L�</&q�N �F�)"|���gX��L��SSc�U5R�7$9!J�=%^��3�b��RE���2�S_�@$�8	�����ư�[��4Ċ��6�T�'�����iȄ����%�� h�࠶i��&:����+�к��������5-=Q�`�a���������?��1��K"8���Ti��)��������x�,�NV��FJ�����Y�>z��-��Ā�𸠘�Ja�$:ڴ�J�NL�	kׂF��)(�ڷ� �O ���/R�:L�G���#$!6F����`��k?maZ�8P��q}��U�|'酸)*-��'���i
��4<������	.�]��:zp�[k�����J��l�4V�.	�`�aٴ���7&���/�>�``�23�3
����}����$�\g�)J$�/��䂊0Cj�5�N1U]W/5�09A! ���F�Q�d����>�׫�l������7ܨar⋿yN��������:���e���2>�R�	��뮗o�k��"�t`O��-Z�"�i)\[�x��+�8�Y�����J�)�0Wj&7�Z=,��0��6RZB�>�7􌍊�MMNn��Meg6*�H�[�N���tR���:L�g��}�/w(�1La�+G{d�g��L�F����^z�e}Y }���mG����S���]��7��A%��c�ڥ+�X�|�E>ߗ#�ۦ�S��$=8[.��By�����\�Q��W�4�7�BX�Iq	*��wq^n˘��V��c��p#��Ȑ�O�\_Q�O�։�u[���E�f`�9h�o|H%�ۚ�%~xm�o�R�� 1qQn��!�i)tL �7��<9�K��)={�ɱ�J9�kp�N8t(�'��9�"]����z�_��v�q��%�e��"Y���2gd?�����6y�����n2ቷ��m�e�����j#(6;8�a%Lc�c��JbZ�N-H�I���j�5E�2}�:B�&ߟ����uyM�]a?z�dF~N�CN�fB?Xެ2������U�C��,C�$,�Z�J�"���0������	xL�;�������S��?�N�{�}���\7j��N�Vb�5��<����[����*�ҿ�l�p�	AQ����*!��r}�K=�Վ,k��Z�R8���$"F�"�=�&&x82������0���{LJ�*�����Q�3D�I|.�5��Y�c��r��1RR�	���g�Jy�i���3!��i��׼��7��w?��L;N>����c���H�K{�����訞��H>8T$[�ʢi$�"O���M��U��%�!S��9E�Z<��=���+9{�I>,���8�E!�(���'�N�X�`�1�PXz�	W3.��5,�ӭ^�Xٸ~yIU�{5�;3�S+7�5����T���}���#\�&-/�S~l#5�<���r�r�T9�g��@�~韒���c����2(�)�i���?����c}����}9��2-7�T����d��R��ۚf#G�d�P�0%!Q�(�8����=zH8�t���?�s-��UVw��!�jT���\{�m*��a34Қ�m�06�c�T,B��5�<��as �շ�jR�FX�9t$G�z�צ���\-D�B�xB���a��U<���: �y��𑹮<!\�>�C�8��!I~���Ɋ�)Q�5�p���GA���hVz\��� �����q�����k\S'"yg|�5��,��h�[�a��2n�(]Ga̍����2i����A޳{�>���2?����ɖ�l����	��Cl�j%�6�J�{�Y�8�Fg��?6<@<\�f�s��c�!֛1Y�:t ���� cE��tAk,dZ+�0vv,?_�ؗ�L�g�s���(�q$'&���63S���(m22T,1~D���4�~�!�au�Sj.�w�29��j���!���9�.+*MB4,�+��э@�<OV:O�D��!b�4�C�UE�r��冨�F�ρ�{�R�gpD���K��k��P9?su��ە�	ۜe. ;%�(�u�%l<�4���L��g��P�y�)5�5�f��=V7:hq��bh5&������)�?��'C���U�TPLǰ.hRC�E�����ӌC��3DO�i9]�Q�Z;*�(��f�Q+���:��\Ņ &8h�X�м�%`�}hZ�X�B�v˼%�N!�Nh�)N��BG�°�rOՈ����f��q!����zg�vD�g�֭A���/�(�᫗�h]�r8�k>�庖��]�Ȑ���4;�k+sg�RyLm�K/(�S'L����[��h�����b~��5�e��,�����̸�~�u�q!�C�i�r�C'W�-5>Ԥ3��h��1��c�6}�Ţ�LU�T���W��'B|�ť��J*��1l���7Pe"�)�°�Fa�}�T?^P 5nOc\�ᙄx�OI�E�j��� f�p{V��S�e����l̥:r�d�^"��g2��n]���u���OԈ+�A6,�����E9L�3B�B��p�����3��3,�BΪ������c&�sIumM)N�S�ݾz�盿��}����=�{��Ԥ$ٶ{�R�������84\��Őz[�QgX!�V֬�B�K��Y������}��L@;����x2�c\k2�d��5�pX�AsQ�p:�-������Gw��5:=b���b�J,$O��j�jӦF��}����N*��Gseߡ��Q�^�P��\�`�&k�FJsX@��	X��kx�%I��QC����KϘ"CQ�pޓ�Pe��zKR���<l(&	?ãb�"+5-z&C�h��b>�̴W&#4��%�a�F��b'`���!��P
��߈/��5�/�k��&�����}o�����T\�q!��M�x��"W��6�Dt #��8�o��b��M5�^4�˄3{�d�������&�
fu���nL����t��}[s��8�rݑ�1�&q����y�<�a.���}9�R��l�A��������5j"��(b���KdY)İ�A�ٰa\�������g�x�й��Y�f/��� �ȫ�c�j9@'4S��\f ؟�-�%�����o0�c��Ο8I�� �{%��%7��عS�N."B��m$�D麜�b�]9��ѧ�d��t�~�����4 "�0�ͣ�Wwbp]GBҵS
�Z)+�Jb\$�89�[.5���T����^B&�\�� }�Ƭ�i= ���B'60J��$����f��V{>�l���+�a�~��+�MϚ&pH�bUX���Z�ǐ�����g�t�(E�P]�5���<��jo��������
h�1i.��	JKp�GO2���Dt��;l`��k5�����\�e�٭�>ǰ��5"#e��-�Rc��3*�}k-F���.:/ѣa=-�y{.�[B�^#gc.��^%X'��. �k�հ���ݾ�d:D��:Y0�нIҽ{���2�n�T}��`qA���w��}��N)�~�͚~�)�%�Z���sz��q���<:ڣ�w�MH�Q��7߰cX�'4Y3��̙39g�3�����+�S���;-k.���`��z9�~���Rвt<��������l;��y�Ms^�%��bť���ﱗk[�K��'D�y=�T�D).���㵒-m3����2��W�c �f�8��tZ�ŧ�5��n�Ϣ��9Yh�L�9��;w���˛yG&�������c$6!Q���G2�o?����{�����)���_r��K%�A�N:W���ǟ�[.9�|�����K�}�tٕ}H�h��O$���?�H��#}�������̸h���-;v4���Q�j�9��T�,���x���f\��϶1�T�2@�f����q-s�"ܺ�ܳc'Y��<��_�,c�{n�����8l��q˭����e`��2������V�9Zn��Fy왧d����E�'��u�˔	�d���d��e3g�5��櫮��c��'�|-�C��ˆ�^�~]�ɂ�W����2.��2Y��Fs}�>9�0�N
���!�b��%	~��AL�L�d��m3���=S�§� �hB�w���-ȕAX;|�����]V�)��{o��&y���M�7���Țg��cǎ��K�� ���C��_��7d�޽�f�RY��q}�9�#�Z)����W��uk% d��+d��G%^��#��Տ��7̞#k�{F��ۧ}����H>�5����B8��+���ǆ�\I�v�pV�`�`z$%3V\�,��~͊<#�X�,���-���9]�Y�?���bhVS�hH�B�C�1��ߣ3�ϼ0�1:w��~B:����.�\�\.#��^���_�X�&=.�P�]-}�t�i�/��-Q�N���,�O���"�o�"9�XU��.Y(�����-�Y���Y?_�TF,�\t�,z|����Y&�� ,],������n�V3 sf
�iH�\���|gnո��m�3�G�չsg��3�r�a�Ŏ���BT������t*��"���y�ҭm{Y��y��7'#����o�U{�i;x��v㍲����w���P�s���ȸ�9��SOȵY�'��,����ˬ�W�ʍ�U|ͼb���目�%��>��"㎛o���%=�w��Y/��̘|�\x�YO�3�-�^��P�GnA�	G&��-��JW��z��L6?#�����-��c�L�ϋ�p��`XĴ��geb 
^1�P+q_�b�n���%D�ʚ�Ke��x�q��ƛ�'6���ǖ,�'�K��ɑG^(K@��0>b��_�<�x�
NYNra���?�R:�ɔ�P�]%1�yf]y����8�~[�L�~�WR
'u����Ҋrs��J�mR����a�r8��ˈ���r���t��bs
?�C��|6�#��a�Ø��4n�rq+kw�9:X�xb����U����b��;j��7@���3��ëW���@ �l��s�%�/��3f������L�`�����!�������Z�r��<�Zٺw�<qw�豺{l��U2�O_9w�D����^:]r�
T��)��� �f
3I��9��z�ϤvF]gaeqq�6��3:�z�I�F�h֢��%�Z}@��B��0p`�^2�����_�sF��8���ԓ��9�\��e x�wʓ/��Ș	�=
N��s��>�D�δ)S!���̋������aw�h�ҭ�����Cǌ���Ζ�O?)C`�>x�=�����W��1��S�,�$?�;@\\����b}��AQ��iT4�~�V7fv��U�so6�`��o�uP���XKq��pY��!)��i��U3f�����ϗe����*Y��?��Nn��P�9),(���Y-iIIҳwoGiIɺ�|!�>�7n�̇eխC'i]�TB\��Ų��/�Uʺ�ou���
Y�{�jj$���V�T3�b��|�@R��T9RX �V�L��VK��/>s�E 0�B�A�J}r6-r��(�Ntv4Ɖ���^8�u����lG�����wh�2
�"�]lb���+.�H<����4b���:M~�|��s҂�qt�us%���9��eӥ��!��\q�����R蕻o�Y�ٱ�.��λ@F�z���0d���4\�uw�� D�W�m��a�_/�:~4O��Α�P��x}���%����#R�9�h�t9��8�6��iA3Ī����|�-�����:ey�2�S�0s���*�.9�<���D� c�e�C���I�G���Y�=��\5�Gk��(��t���?��};'M�U��W^�%2�>���INO����\��J�(+�?�q�m��/�(��?�q���i���uS�W�LO�zNyy���U�0����U�@\���2�
�e�v���5}�LE�&< 	��1~�Іw�63��*Nkiƌ��:����RXX$� ��S�X t9��HO��FY��S��8b�P�鐙)�m��#��I8f�������D ����>��Yet�]��4^����Rn�s���\1�إ��fΈ桅4��N3�[�f�5'a�-�{ '�!옙Q�$��"���y�I�K��
l�D4�?���,�������k[��-ǎ�~#I� �#֩u4ܱ ��. �&���Y.��'��Y +k.y*��~��r^��d���䣯��E8��w˾�#�ze����(� ������;}y��3�&�F�q�u�]!����u�˒��/�l�/��#X�$��N#�-u���+N�e�z����OL��HԏG��$+V���n��u~I�U@�k���\�	������`P�{}�_� ��	�_t1���r,��z)E?x�Ϥ3�������/a�>
�롟�)�m�{O�b.,/�m�w��{�W����o������-[���q���ڙ%��t�t��C���q�{�����b�/���'�|�Y�Z1i�V��J�+�������r|��2+�JW$�3V�x��Y��l�^�LE�ڗ�[�0"�]z�&�);��� ��}Ë��(XD�ګh��Q� ����iBg��CK�{�"��m��{�K>x쨼���э�5 � t;XE�u^y�/ʐ~�eǾ����oj)Wt�����^X�����]Jn{���U1N��t�B8X��)E��U�i�a�N;�h��G��'g՗�2H�)h�ְZy���J>	�ʰy��eݳO�m�f�
s�c�wΙ����g��k�]*�;u�����o��Jy��Wd)D��5�{\u��Ɇ矓_�����k��Y��C������?��:�'�>����	\���_��q[����4pnYA�Վ�H�����.��2W�l�@��bs��~V-*RE��#Q�:`e�4���"i�Y��\��-�_ Q)�V��뮹F,����*膻�ܠ����K.S��{o�EcSD��y���Bde�{��w��?���ҹ[W��?>�5�{��W�����X�>����3�T�E���"[���D�iv:5�T��|���J�.	"�����v-�u�K��ʙng��	&4 ��d���e�!�kΚ����b�&!�3�`�7�5��Æ�J�*X>]�w���V�ұKgY�B]Go�!w�^2�f�XS�:u/8�Y �e0�6������ON�g��+ŕ��k��ևN]���c�>2t��:��hMZ�ԓJT渃������k�B�/��8�nۧhL�kYP�1�����O�b��BM��î۟�6r�R�����^!w���Y�z������t����@'7P�R�ρ����3��%��,�/;.!�he}���0�_��8�LV���G��d��zV����'����A7v.û��E1��\�͎��%D��V�l ,����T��(de5��C'u#���#�e7�����f;~ٜV�6/>W=�y3I�ef$�X��+'_,WL���՝S�A�����Kgmù�/��By��7e��ź=�� ��/��`���!K�u�*�߽��,��~I�HSK��Kuiv��]��nVq�=<�?u�r�G��\�����҄t.Q@�s�nkr�}d�~�$�K(��?-�'b��&{0(�2RR5�S��L`�Z�"�8SA�|�#,XaYY�����xS�d�ȊpSS@�k5��k����)�)(�@dw��"��/@uj�^�2ZP��Y�&��o�H񡼣��o��tTz��6��={j�q��*}^y�4�'�ڬ�5�M�
�j+"�g��یz�<\9�d��`���u�Zv�">��.)���)JU����55C*�m�7G�L�S�����g��Qce�E��?�~�M`�2�y�5b�)#E_瑊��t�5��:y�����#��v(W�5��%e����J⋯�Z�G�X[�>o�1S�OhP1a��B�yh�|��7 �aE{͌�r����ҾM �[Y�@������V<*��L�	�����V�H�L�d���Jp4C�p0k��8�['A�9|X�⫪����_%� ~���콠�5y�MZX��s2ȸh�E˺�k����o@Ɯkg�J"�1n�x��O���dpĮ?��	�z(��Q���@��Y��s�\G��ʫe2D�$2n�3G6����;�[￧k��7�u�fF��
JJe@�X	ۻ �y�6@t��-?�Q����'���6NL�'Эc-�싖[����;e�͟b��� Lsì�$��&��{��g%?/_f]>]�)����g��eM^�aT�R{C�S�����c��3SӤS�.p���xi���\b�����N��$�ظNk�N�s���u�GA�U��hp�\�a���'�.z�iu����\wx��V�MsMO�1!@j�D���YŜ#˻?��`�Gi~�q3�q�1�X�!iY�!v�=��%vy���l�&h۹�D�½Y(�9Z�������V�~�-;��;XN;�ee�,u�[�>�����M�[��ZҦ���T�P�Aj��,{K��P����43�Z�ݢc�a�יA��������[2,��;v��3��}�޲�LC�D���]��ܠ����N�NIL�^=z4fϋ4��`8���szë���&��υ�����3\H��\;�R6�Z?��۴"$����� J��Zqr�^��4~+��r69�}zI5 ӹSG�ݥ�Y��k�����7KdF��;S=m��9�{M�+�Z�P�rp~ƔiR]Z�[����ʆ�s/yq�q�רes!�6�X)����GA��{���'��ku��P�E��Z�oʔ)Mr���յc�.�b�������A��C�s���r6���i�5zA1�Z`� e�;-�lw�?�	X�2�
�	�v<���t���l%L]��e�x�cm͹%"G,#�"����3����r킵I(D+Mm�q��X�J��-O�;��++��:����3L�a�-w�j�Ch�Atf[��1���6��`�(�䶷O3F6>�Z��Xٝ��'=�89��ه�ް��*	v6{wp�ry��ݽDH�Z�͑��o����L��lBІV]59�����uVM�{�]�����xʽ�h���9�g��[���E�9�f�a���f�:�c�	9�U?[Y�4[Wwb��6��Y���[�Ĳ�dA~��ܹS�!:��)�*&�##��!Ԭ�ҘO�l�P��İ�]-�2a��ս��$%)י�@����Y�i����V�]�����ʎG��I�Z��v�M��ptę+��m�t�Kp�[�!6PN����;Ԇ�ݯ��W�����p�l �}`*r�rR!���wLJ 6�qh�}X5�l3V�2��Yج�*h�f%F��'��fp����ڛ����zS&��{�}a��W�$6Nu�g�<ے�K�US�"��Bq��.�2��%�X������Ĭ�ON�F�_��ע����!�f��i��f�?�bW�qY?a�<�>+���a��S-��P�!h���ٕ���C�ɷ[�4��T�v	�.�9�[��(V�{!Fs`��F���ڮU�Y� ��r����Y�{��z~䐡��o�@�ڹ���UD&�M=F�ee��h���f�6�C�4������u51���GU��g�:g��ߏ�+��=�U�Ox�k#��4UTW�����}�NS��;��:�̰�wRlff��O��[��mI`ۥ��t3������h����Me�iJ,�8�W!�9��;�Lnjav�8�q�Z��쵌`����6�l��n�^���qܧ��d��]�T��_��Ajj ̚*M��=d�I\M7�;C�5eFx����~��}P��q���={�xL������a��u�u�&����ߟ|"Eǎ��d�4�sss����-�4`��m�n�vZ����D  ~���p;L�)cA�gζ��uK�qWTʷ_%�� �u�!�LZ����	׸t�r4�<�j������ښ�j���KL��/�kN��qKC�8�M8�c]�G'�aL�� ��Aݘ��-���o��R�yM����&�`C�E67��-T���VM�c���G�g����ݧ�m��⼜\1i��"ɇ(i����/���@������B����TfBDr97�1QM(�ҍ���꫔��X���dx�㡸K��K�H�;X,�32�@��ȑ�bIOMwR�f�Y���V���zt�̮�σ�;�������N��f�I>�ݠ��(eg��fE��H9�S�ԟ�%UU>�*o��P�п��dae�Y笠M 0F���v�̝��}("���W*��P���QT����AZ�$�a`� �m�OSbs��ʆ������=�|o��9�V����9����B����n����$�F��3"�&jw�CM���C�g��q���=~��H��V:Y4�d���2�\��5+���ū���[arY���~���L��k�w��Y�u몲�:p̘�z/�l��/8�|��D���͝_����9g�~g?�:uԾt#�a�飐"8��~}�6�C�bҤ�����:u�ϒ�F�a����-+���N�oP��{pl���&yYg�.k��q<��0�1'1#�a�eɉÇ��ޮzLz��ۆ�m����r�u�V	��aV6u9V~/�
~��\��qj�e�kLFs���Zw����F��\v?a3$�<|'�\�-k��n��q�?:�.��O3����aIB?�☋#�,��|4컩�fk��o{�BTăb���P�Bv�!y�����(�k�;��F�c��*V�޺Vv�T�4��V��LZ�R�~Z}g�5	�G�}�g8���� �L��%    IEND�B`�PK   ��-Z����U  �  +   images/e1729bf1-0a9a-41a3-ae0c-c5916288453e��gPܷ�C��(U�HQ�5�"RC"��T�
�_D��B	�J�.��zKB	�����9_�{�מY3k��~f�̏�����X�@@CCx�� � N�?�3���������C� �a�����������������������������$��@��p����S'&1o���>~a�~����l'���'����������ԍ����UT��<���d�����
dmc�����k7w_?��������ظ��	i�22�>g�|-*.�V����G�����������?�spbrjzf����Y][�����N��g4 :��������CKOOG��ׇ�6���<�eS&'�+bw�1s������庂����8+��"Z�W�?F�wB��_F�+��>�y@��W��������/�D����^f6ffVf&&���l�`b��q�������ߍ?�������	`����m�8@ I��@D��§ۮ� ������ٲN�CC����;E
�P�Q5�Ȯ~�3$�vo�
-25�PP�����X�Τ�w}
3	}	$�܎'i,=���%�+��4f�Ԏ[���t�Difkf�~�� P��`��[ qY6a"^ۗ{��)j�[��)�B����|F��v�`�c�Y�n��m	dL���5���E��I�Y������fQC����k�K-(��y��
����7�V#����:j���T"4��=�&J!�_9j�HJ��.���
�}Aۥε`��~lk�b�l�#�luv�ڳt�o�����u��L�P�#_aЩ=`�M�1*��v�ػ�:�q���3�h���C������&��vH�!����b`U����N�&����7��f�,(F��z��"	���r�pp�'�}nH�a$�;�L�Mw���r�v�����1�kG��'=�T����E� RXu&��۠d�>,�ѻb�
Be��/LR���'R~��Y�~��=�����<��i� �*��|(p=�Uw�)��"r����I��(J��ُޒ�ʚ�����'�a�`�����XS����\�&g�˰�i�*;�P-��F���oy�dM,�O*��(�
��$7Ԯl�;�]�;���D��N�v	l"������n�O"��^�����9���L�K���W��6�<���[Bf�t��L�m�%�6�sS� ��2�(��-n=,ʛ�0�J�� �
�:R���?/ǴI8>��I+��'�$��Q�U�^醂&
ܒ�W�9�{GtG}�o�9���/�Pn�0���M7
�/����2'$I�T��@�+����#x����w���
�OЛ�J������?��/�����y����@6#Z�:�/K�ثA/�&�Zй����m��o>^)H*=�m7��<����W<]�[mg{'{����s_�%9�Jv��V)׺�����M��y9�}�ȫf�Q�}J�G7��ubнr=C�
���U���e��D�>�X
���D����~a�M	#"='>��?�t�N�^= ����:^�:e�x�e��j�+�Q�K���y)�'��b�jń�ܐ#9���h�b�ձ��V����g� S�֚�St���l�(��ُ6�Ý�+��4�E�?���ҵ1���3�:�)�1OM0%?h��**_���]�R����FI��b��_��4�c�Myy�6�{��|s1��iD�J�k������S~�gsC�
���6�ε4�EU��x* ����&�nG���P6���/c���ch آCF�~��w��s3���G�	g��nփ�GNE���?��Ңg��s���փJ�T0c�T 7�ƞQ�}�6H�J̊NI��C7���sQx�� cw�R�є&h�Юd���գA��]`����oW��-�.�Q�8��6�)�>�c��Ά}��L�u�^],a�3�)n|Q�]M��duZ[p�"�/�'_)sG��S�f�Nͭ��{6�j��GѝjדjF�	�E&󻥨��@�]�n��2�𪀝�ߛ%�:�ҭ��H��s}4.��0�Ē��>z��?���V;(��Lc��9���6?�rNƮ�Qd�:�ɳ�5C��	*�\8��2��C�Se�XP���6�
����7"�W�d%_�#)�S�7-_02�r�^֔P��P�F"����2�9{�
��5aO*�yDA&������k����G_�`�i%3|�5�������a��`?�#>��C���"�S	��:��a͈d��oB!����j�2>�k����������/����,�y���f���^m��r��u��0��N~g�)��|+���Al���'v�Ei���ʯ��MB����GAa��5f�_�`��y�ԅ�M�����XE���b�8�NY�t�7��>t���bb>���a�=���*�FYE�;�7�#����vo}B��O��}*��@Q�O��c�i����T2'`�6K0�c<4�����uʃ)	3�X�P�"��?"�3���p�l�R� #��=�7~N��鎲�o�@�!5��E�CǮ�� �e*ൣ�.t�J���g�+Jl�˪������~�qԚ�]��h��Zś�`���T�&�bz]b��r!>NeXS�Iӄ��Q��s�HEr�]�:����k���
���{U����~�eK�k��6d�H�1���w��	�xt�]O�W�f_]߻�[���;-��z�N�
�jY���ȩ9� \�Y�y
�����Nի����6�~$vQ�B�(g�*2�bI'	Āc�$�������׶���\B�^��۴y�cJ$-ã4�I�7�Y`Ę�eA�Hu-x���	�L���2���z�qK1x�~�0��P9�.�v���e�>t5r��6��-*eQ-���|��OnD�M�-��Yl�gzv;�Q�+�Q�)�_�<�����\)v�i@�3���U�4]���; /z|a��3��J��Pl~���o����iS	��9�)J�kh����.��C��x9�p�!R��vE�3�[�+�Ҕ�ثv�1���7�0���N�>ۤ���+���:���buP��r�?�s��F5��`�~?���I<}:�i�!��\G;��35��.��o�b��{��������?�AAW��1xh�D<O���۵�c���wǃDH;�;h�$����9,C�_>�p��U&�Z�}P�uS� V��P:�U=��q�<�����ќ9�گ��Ȱ]���Nm�|��m��O����VK���t�$�'VZw/����T��f��K�gy�.zd����W>��v�Q�$��5N�+�3�C��2��J��YD��ǧ@E��@f*��(A�kz�{�����MP��Kᚺ~Ot����7�1>��J(6g`��[#ͩv6��9МK/�uYo��N)*���m�YͿ�M.��c��#�v�üޑ��M�ZP_���y�Us~�(	���&)/ľ�qG��9ϥ7�{%"y$�Z�x�a2�ov?�^���~�����W��y��~c�M@.�����<��͋B�~yY�u�5�W|3�<*�c�gG5j/�K���3�o��Y�I�G#�?��əæ�`�z�>krBS{Y��.�b�}�����7���ߘ*�L01
��l��u����I����Nb��~}��3�c�
��'�	��b���0����S*�z����M���L�4EJwq�Fz�w3����mKb4]c& =�`��W�o���dGB
���*�o���̩�([��4��<���Ѡ���C9&��Wr���uEA�D��o�H�4��:�8�}��쇓����5�pY�c��%,�t�`til-|Q3U�� Ϫ)}�F%�{Y���[&���!�`T{��or��B�"��o�������Ύ��m|�	|�>�?�	(���ۤ�De8@,�e��o)H�H�<��G�1�����Kk��;1]z�Y�'Q��Vi�۷�D�a;4OV&Q?�/�8�W�-�4���NK�^ŔNA�x������Tb��[��"WS?��&	~�����xv��e�e��0$:LeP����[:ש�C���I���Eu��S���Y�Η_A�>��)M��KAQ�[+��J-����i68�b���of�D�T6�;K��K���#[ ��:~3��޻҇���m��>���u�/����7��ZǪB�5	����k�-�fK���\e�0�s+{�.��kR��d����
^�\S^؆���I�T2#bg��}z����^�.�R��A�Ǒ�K�x�&�z�ʢ�ْش���W����O�Y|��i�=�{ʣ|2�����_�Ӱ�<��k� lg�'�(��j�����ۥ��ݺ#}
K�ǹoD�R�0����N:�R8!ßDN�/qWa�&&����j(�=?t�W�ޮpH.�a�Hj�X[��_Q��o�7w��F���'�vڂ��o����,����݊�7�x���n���~7#�RG�P������o��
�_+������!�vA�����n�?�M����7��Vő���'��;��?���'���[��F�D��_Z>K�@V5��Ŀ0��Ǘ׿�B�U���NO&`�!r��2�܏kZ����G�����b�	q$�⒮r�f}�ە]�fX}lQy�H��]��S�<HI�Eo���"˱�R��zl\���XK�����&��*���;*�
ȇpC���BL"���Ҷ�R�������b�O��n��	V<O�P��"��A�]K����5��uf�&���(6W7��c�\�<�����v�����������������������f���-�n���oF�K�˷��5Յ�?r��Y��`�m�z+rXG�^��F��_>~v����F��d�s��ܕ�yP36����\�=��g�J�������g�eX���(��'[䉎N�9��u��Hz��X�q����I>�w~������-��Ů�tj��FI�.�"���M$��tI���%G��7���v�{��'")�ObzgV�_O�����Q"�	|�'��Vr� ,�#�S� ��rT'�h��O�-*���6Հ�~;ctm��(\50A'$�w"��&L<^�P�������(s�����1�!މ���z;���9�wM~C����q�WӒ�	�F��K�p�T�wU8�%W����A�|����}c��EY礯o�X=��7!��8}�R�s���!"`�s<{����29�V��h����_��m�  T�?��R�/`�;�ٰm|��b�>N��]A��#;�bpg���t��1�O��v�B�F�e�
��κ,ṃ���La^tV��_v���:��)�P���V@9�c	���9�O��4��aΔ5���[�e6��"���f^�e�G��f�K+@�=( ��9֮���L��[+%����"��T�|"�N�B����#-I��~�=Nɋz:)�X��_����~&�v���c;7I��Nv�x��pN|���Mx���bA	��n��X���(���R� W2��*��"+кY�T �ݒ������Tqt_�Z�W=��Rraf��{o��;�/���$��o���<l��K'�gy�jX��w���ois��*�r�b]$<l�O�(S�W4HAE]!�-+�K����F�N+�
RX��U4�O��s�I�/I_�Tv��{`�
� ό�K�e��ן�������fdm����|�`�T���<	E1~�idl�Qh=�C�eL��S��=SG*���X�������"?��R}T�e�ʠ��F �x�A/+�����n��T~�x��g�II@X! �B�5�J«�Dm%Y8�����pq���s�8"���g|���T`����A�B��ba�W��:���&��x[�dΨ���)��Sm����=��J����Mr��iD�_�"�F۟�PR����Fߺ�2��U�yD��3م�\1ً=>f)Z?#q^%��A��k���`O�ႌ6��C�7d�����H���A�j���n�E�x��PP͊[�
b��n~���@��6DZ��)�c���n�#4�:�O�&��������?:�s�㝎Bܛ���X�v�^��c����/|�|Q�	~@�l�P��:��Sl��S�Ze|[���xL��!���qT
�L!נ���(�2��kZ@')� 4j7�H�8_����;��-��5���*�ť��6��-M���7��T@V&\�m��׺W	���.�P�x���*`~�w,Sn���Ӎ�Bw�]QJ��8rN-�}�
HV�lY�1���a�nl�R5��wy��O�"��hWMP��"�]��B��o��a�{�6��*�[=�*EC����M�P�5�}K!u� PK   �-Z��:�  �"     jsons/user_defined.json��ko�6����}� K�U$�-s��XI�v����V�#��ݬ+��G];��T� lY<y������t�e��g��F5�sU��ʧ��g�lʺ�?��P?��������ϯ�/��m{�仲�'�/��k2yS>/u�LnՇ������O_�YSgu�m��J5�w�}1�϶�Nͦ��4%y��"gy�,GQ��rJR 2�8��]�M֔�m����2�߹y��4"Di[2�� ��LeLr��u�A�+>���w��Q���������r_���e���zz�uZ��.��z%���v���!́~���u}��b!!��ޝ�����=��Ͷ)u7����M��e��OX�ĺ��3!����rs^e�F7�;o%Sվ�|�|�mf�뼷N��z!W�#�^^8�#ük�����i�#�u� 3
H�0�a����7�N
�R�! 0�rq�P/��0�NQ�-v A(� �f����0ې�-N�ˉ^.7WlI�Hp2����!���S�T�����@A����bQ��W�(�eM�yk��)��!Ա�#�K�X��r��M0e�@�������'ښ��E�D#���<��T9$cG�"�T9� 	�[�}S�z�[�H��j�T7d�' �↼�e�B��K7��5������LE#8�����!Y�m4ھ;�!ˆ=Ȍ�`�n	 �VM����w�:d٩�h��mߔ0�>������8�L1 �!�$��j��;gB���)���S[�|q�t瘦�Q�2t� ���l�����j�fX4}���'pc�������|���H�<~�X�}��w���"`8���E��	w���v�p�;Na�N-�Tc!q��[u8��	��!� �N��	�M0��O��	�M����s��s�Ē|�� �Y�%�OA�eM,�7�C��[�Ē~���vD,8�p��w"��ŀ1�r�)m�����,��+ѽ���e�rM���z��mٕB�+eVW}�QR�s�Y���#D	BQ��,#��c1�;�A��39�+W���}&���-��w�R��v_���pW]��ݝ~�J�/r���}Uu]_V�%$E��BD9LID�Q)	f	EhYUp$�,ǑR,�t�,�J���4�E��ȇ?��^u�ϡȹ�M���{�����LW�p��}�z�O�lZ}��r�k�l���IZ�=�1�w�V����ɶ��������+hۏ�Q�v�wU������'������c}��tw��l}6-V�z��e��7���Ճ#�FG]8�S�����wU>�Wus4��wac�\�e�hPp����F�@�7�WE]mo��Qg�Lud^�R5�Ku���#=�4IrP�
��I�+���8d� 
@��au���~��z^�2֝0���Z�x���A���A"AQ!��34�$U0������d�l	RzE*�L�-S����E�@*' ���S�!�0RȈ@�u�E0ѹ(�X���K����2.Y�~yɂ �Y�T��h�Do�s�⭙��������t�r�}����o�Q�,�Ą� S������~�q��i�����!��0Ƭ'��ӄ�|)��HqZ��B1
������G\�V�<�~:	x�Xt1l]?�RZ��c��V#���A	�s0�s��N�0� xNr���r�bg��	���gQ�=
�벛��,&��9M[nP��O�,m��I�<74?�_�,�4��'���c$F��ܖY����"�?'.glE��8
��q��}ĵܝ�rӐ%�>�[�N��?\Dcbܛ�˰3շw��PK
   �-Z����  R�                   cirkitFile.jsonPK
   �-Z����7  �  /             8  images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   ��-Zl��B�  +             �   images/60459fb9-c9d0-40e2-ae43-752ef2ed40d9PK
   9�-ZE�U� z� /             �" images/8a9df60b-44ed-4a65-94c8-aaba687a6de8.pngPK
   �-Z�&�}[  y`  /             I� images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   9�-ZG��{p5  k5  /              images/a528d487-389d-409b-9452-c3cc4275f339.pngPK
   ��-Z����U  �  +             �S images/e1729bf1-0a9a-41a3-ae0c-c5916288453ePK
   �-Z��:�  �"               nm jsons/user_defined.jsonPK      �  �t   